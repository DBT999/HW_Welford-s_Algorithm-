module inv_x_count_LUT_prev_and_next #(
  parameter int unsigned
  SIZE_X = 1024,
  WD_REAL = 16
)
(
  input [9:0] x_count,
  output logic [15:0] inv_x_count,
  output logic [15:0] inv_x_count_prev
//  output logic [15:0] inv_x_count_next
);

  always_comb begin
    case (x_count)
      10'd2: inv_x_count = 16'b1000000000000000; // 1/2 = 0.5000000000
      10'd3: inv_x_count = 16'b0101010101010101; // 1/3 = 0.3333333333
      10'd4: inv_x_count = 16'b0100000000000000; // 1/4 = 0.2500000000
      10'd5: inv_x_count = 16'b0011001100110011; // 1/5 = 0.2000000000
      10'd6: inv_x_count = 16'b0010101010101011; // 1/6 = 0.1666666667
      10'd7: inv_x_count = 16'b0010010010010010; // 1/7 = 0.1428571429
      10'd8: inv_x_count = 16'b0010000000000000; // 1/8 = 0.1250000000
      10'd9: inv_x_count = 16'b0001110001110010; // 1/9 = 0.1111111111
      10'd10: inv_x_count = 16'b0001100110011010; // 1/10 = 0.1000000000
      10'd11: inv_x_count = 16'b0001011101000110; // 1/11 = 0.0909090909
      10'd12: inv_x_count = 16'b0001010101010101; // 1/12 = 0.0833333333
      10'd13: inv_x_count = 16'b0001001110110001; // 1/13 = 0.0769230769
      10'd14: inv_x_count = 16'b0001001001001001; // 1/14 = 0.0714285714
      10'd15: inv_x_count = 16'b0001000100010001; // 1/15 = 0.0666666667
      10'd16: inv_x_count = 16'b0001000000000000; // 1/16 = 0.0625000000
      10'd17: inv_x_count = 16'b0000111100001111; // 1/17 = 0.0588235294
      10'd18: inv_x_count = 16'b0000111000111001; // 1/18 = 0.0555555556
      10'd19: inv_x_count = 16'b0000110101111001; // 1/19 = 0.0526315789
      10'd20: inv_x_count = 16'b0000110011001101; // 1/20 = 0.0500000000
      10'd21: inv_x_count = 16'b0000110000110001; // 1/21 = 0.0476190476
      10'd22: inv_x_count = 16'b0000101110100011; // 1/22 = 0.0454545455
      10'd23: inv_x_count = 16'b0000101100100001; // 1/23 = 0.0434782609
      10'd24: inv_x_count = 16'b0000101010101011; // 1/24 = 0.0416666667
      10'd25: inv_x_count = 16'b0000101000111101; // 1/25 = 0.0400000000
      10'd26: inv_x_count = 16'b0000100111011001; // 1/26 = 0.0384615385
      10'd27: inv_x_count = 16'b0000100101111011; // 1/27 = 0.0370370370
      10'd28: inv_x_count = 16'b0000100100100101; // 1/28 = 0.0357142857
      10'd29: inv_x_count = 16'b0000100011010100; // 1/29 = 0.0344827586
      10'd30: inv_x_count = 16'b0000100010001001; // 1/30 = 0.0333333333
      10'd31: inv_x_count = 16'b0000100001000010; // 1/31 = 0.0322580645
      10'd32: inv_x_count = 16'b0000100000000000; // 1/32 = 0.0312500000
      10'd33: inv_x_count = 16'b0000011111000010; // 1/33 = 0.0303030303
      10'd34: inv_x_count = 16'b0000011110001000; // 1/34 = 0.0294117647
      10'd35: inv_x_count = 16'b0000011101010000; // 1/35 = 0.0285714286
      10'd36: inv_x_count = 16'b0000011100011100; // 1/36 = 0.0277777778
      10'd37: inv_x_count = 16'b0000011011101011; // 1/37 = 0.0270270270
      10'd38: inv_x_count = 16'b0000011010111101; // 1/38 = 0.0263157895
      10'd39: inv_x_count = 16'b0000011010010000; // 1/39 = 0.0256410256
      10'd40: inv_x_count = 16'b0000011001100110; // 1/40 = 0.0250000000
      10'd41: inv_x_count = 16'b0000011000111110; // 1/41 = 0.0243902439
      10'd42: inv_x_count = 16'b0000011000011000; // 1/42 = 0.0238095238
      10'd43: inv_x_count = 16'b0000010111110100; // 1/43 = 0.0232558140
      10'd44: inv_x_count = 16'b0000010111010001; // 1/44 = 0.0227272727
      10'd45: inv_x_count = 16'b0000010110110000; // 1/45 = 0.0222222222
      10'd46: inv_x_count = 16'b0000010110010001; // 1/46 = 0.0217391304
      10'd47: inv_x_count = 16'b0000010101110010; // 1/47 = 0.0212765957
      10'd48: inv_x_count = 16'b0000010101010101; // 1/48 = 0.0208333333
      10'd49: inv_x_count = 16'b0000010100111001; // 1/49 = 0.0204081633
      10'd50: inv_x_count = 16'b0000010100011111; // 1/50 = 0.0200000000
      10'd51: inv_x_count = 16'b0000010100000101; // 1/51 = 0.0196078431
      10'd52: inv_x_count = 16'b0000010011101100; // 1/52 = 0.0192307692
      10'd53: inv_x_count = 16'b0000010011010101; // 1/53 = 0.0188679245
      10'd54: inv_x_count = 16'b0000010010111110; // 1/54 = 0.0185185185
      10'd55: inv_x_count = 16'b0000010010101000; // 1/55 = 0.0181818182
      10'd56: inv_x_count = 16'b0000010010010010; // 1/56 = 0.0178571429
      10'd57: inv_x_count = 16'b0000010001111110; // 1/57 = 0.0175438596
      10'd58: inv_x_count = 16'b0000010001101010; // 1/58 = 0.0172413793
      10'd59: inv_x_count = 16'b0000010001010111; // 1/59 = 0.0169491525
      10'd60: inv_x_count = 16'b0000010001000100; // 1/60 = 0.0166666667
      10'd61: inv_x_count = 16'b0000010000110010; // 1/61 = 0.0163934426
      10'd62: inv_x_count = 16'b0000010000100001; // 1/62 = 0.0161290323
      10'd63: inv_x_count = 16'b0000010000010000; // 1/63 = 0.0158730159
      10'd64: inv_x_count = 16'b0000010000000000; // 1/64 = 0.0156250000
      10'd65: inv_x_count = 16'b0000001111110000; // 1/65 = 0.0153846154
      10'd66: inv_x_count = 16'b0000001111100001; // 1/66 = 0.0151515152
      10'd67: inv_x_count = 16'b0000001111010010; // 1/67 = 0.0149253731
      10'd68: inv_x_count = 16'b0000001111000100; // 1/68 = 0.0147058824
      10'd69: inv_x_count = 16'b0000001110110110; // 1/69 = 0.0144927536
      10'd70: inv_x_count = 16'b0000001110101000; // 1/70 = 0.0142857143
      10'd71: inv_x_count = 16'b0000001110011011; // 1/71 = 0.0140845070
      10'd72: inv_x_count = 16'b0000001110001110; // 1/72 = 0.0138888889
      10'd73: inv_x_count = 16'b0000001110000010; // 1/73 = 0.0136986301
      10'd74: inv_x_count = 16'b0000001101110110; // 1/74 = 0.0135135135
      10'd75: inv_x_count = 16'b0000001101101010; // 1/75 = 0.0133333333
      10'd76: inv_x_count = 16'b0000001101011110; // 1/76 = 0.0131578947
      10'd77: inv_x_count = 16'b0000001101010011; // 1/77 = 0.0129870130
      10'd78: inv_x_count = 16'b0000001101001000; // 1/78 = 0.0128205128
      10'd79: inv_x_count = 16'b0000001100111110; // 1/79 = 0.0126582278
      10'd80: inv_x_count = 16'b0000001100110011; // 1/80 = 0.0125000000
      10'd81: inv_x_count = 16'b0000001100101001; // 1/81 = 0.0123456790
      10'd82: inv_x_count = 16'b0000001100011111; // 1/82 = 0.0121951220
      10'd83: inv_x_count = 16'b0000001100010110; // 1/83 = 0.0120481928
      10'd84: inv_x_count = 16'b0000001100001100; // 1/84 = 0.0119047619
      10'd85: inv_x_count = 16'b0000001100000011; // 1/85 = 0.0117647059
      10'd86: inv_x_count = 16'b0000001011111010; // 1/86 = 0.0116279070
      10'd87: inv_x_count = 16'b0000001011110001; // 1/87 = 0.0114942529
      10'd88: inv_x_count = 16'b0000001011101001; // 1/88 = 0.0113636364
      10'd89: inv_x_count = 16'b0000001011100000; // 1/89 = 0.0112359551
      10'd90: inv_x_count = 16'b0000001011011000; // 1/90 = 0.0111111111
      10'd91: inv_x_count = 16'b0000001011010000; // 1/91 = 0.0109890110
      10'd92: inv_x_count = 16'b0000001011001000; // 1/92 = 0.0108695652
      10'd93: inv_x_count = 16'b0000001011000001; // 1/93 = 0.0107526882
      10'd94: inv_x_count = 16'b0000001010111001; // 1/94 = 0.0106382979
      10'd95: inv_x_count = 16'b0000001010110010; // 1/95 = 0.0105263158
      10'd96: inv_x_count = 16'b0000001010101011; // 1/96 = 0.0104166667
      10'd97: inv_x_count = 16'b0000001010100100; // 1/97 = 0.0103092784
      10'd98: inv_x_count = 16'b0000001010011101; // 1/98 = 0.0102040816
      10'd99: inv_x_count = 16'b0000001010010110; // 1/99 = 0.0101010101
      10'd100: inv_x_count = 16'b0000001010001111; // 1/100 = 0.0100000000
      10'd101: inv_x_count = 16'b0000001010001001; // 1/101 = 0.0099009901
      10'd102: inv_x_count = 16'b0000001010000011; // 1/102 = 0.0098039216
      10'd103: inv_x_count = 16'b0000001001111100; // 1/103 = 0.0097087379
      10'd104: inv_x_count = 16'b0000001001110110; // 1/104 = 0.0096153846
      10'd105: inv_x_count = 16'b0000001001110000; // 1/105 = 0.0095238095
      10'd106: inv_x_count = 16'b0000001001101010; // 1/106 = 0.0094339623
      10'd107: inv_x_count = 16'b0000001001100100; // 1/107 = 0.0093457944
      10'd108: inv_x_count = 16'b0000001001011111; // 1/108 = 0.0092592593
      10'd109: inv_x_count = 16'b0000001001011001; // 1/109 = 0.0091743119
      10'd110: inv_x_count = 16'b0000001001010100; // 1/110 = 0.0090909091
      10'd111: inv_x_count = 16'b0000001001001110; // 1/111 = 0.0090090090
      10'd112: inv_x_count = 16'b0000001001001001; // 1/112 = 0.0089285714
      10'd113: inv_x_count = 16'b0000001001000100; // 1/113 = 0.0088495575
      10'd114: inv_x_count = 16'b0000001000111111; // 1/114 = 0.0087719298
      10'd115: inv_x_count = 16'b0000001000111010; // 1/115 = 0.0086956522
      10'd116: inv_x_count = 16'b0000001000110101; // 1/116 = 0.0086206897
      10'd117: inv_x_count = 16'b0000001000110000; // 1/117 = 0.0085470085
      10'd118: inv_x_count = 16'b0000001000101011; // 1/118 = 0.0084745763
      10'd119: inv_x_count = 16'b0000001000100111; // 1/119 = 0.0084033613
      10'd120: inv_x_count = 16'b0000001000100010; // 1/120 = 0.0083333333
      10'd121: inv_x_count = 16'b0000001000011110; // 1/121 = 0.0082644628
      10'd122: inv_x_count = 16'b0000001000011001; // 1/122 = 0.0081967213
      10'd123: inv_x_count = 16'b0000001000010101; // 1/123 = 0.0081300813
      10'd124: inv_x_count = 16'b0000001000010001; // 1/124 = 0.0080645161
      10'd125: inv_x_count = 16'b0000001000001100; // 1/125 = 0.0080000000
      10'd126: inv_x_count = 16'b0000001000001000; // 1/126 = 0.0079365079
      10'd127: inv_x_count = 16'b0000001000000100; // 1/127 = 0.0078740157
      10'd128: inv_x_count = 16'b0000001000000000; // 1/128 = 0.0078125000
      10'd129: inv_x_count = 16'b0000000111111100; // 1/129 = 0.0077519380
      10'd130: inv_x_count = 16'b0000000111111000; // 1/130 = 0.0076923077
      10'd131: inv_x_count = 16'b0000000111110100; // 1/131 = 0.0076335878
      10'd132: inv_x_count = 16'b0000000111110000; // 1/132 = 0.0075757576
      10'd133: inv_x_count = 16'b0000000111101101; // 1/133 = 0.0075187970
      10'd134: inv_x_count = 16'b0000000111101001; // 1/134 = 0.0074626866
      10'd135: inv_x_count = 16'b0000000111100101; // 1/135 = 0.0074074074
      10'd136: inv_x_count = 16'b0000000111100010; // 1/136 = 0.0073529412
      10'd137: inv_x_count = 16'b0000000111011110; // 1/137 = 0.0072992701
      10'd138: inv_x_count = 16'b0000000111011011; // 1/138 = 0.0072463768
      10'd139: inv_x_count = 16'b0000000111010111; // 1/139 = 0.0071942446
      10'd140: inv_x_count = 16'b0000000111010100; // 1/140 = 0.0071428571
      10'd141: inv_x_count = 16'b0000000111010001; // 1/141 = 0.0070921986
      10'd142: inv_x_count = 16'b0000000111001110; // 1/142 = 0.0070422535
      10'd143: inv_x_count = 16'b0000000111001010; // 1/143 = 0.0069930070
      10'd144: inv_x_count = 16'b0000000111000111; // 1/144 = 0.0069444444
      10'd145: inv_x_count = 16'b0000000111000100; // 1/145 = 0.0068965517
      10'd146: inv_x_count = 16'b0000000111000001; // 1/146 = 0.0068493151
      10'd147: inv_x_count = 16'b0000000110111110; // 1/147 = 0.0068027211
      10'd148: inv_x_count = 16'b0000000110111011; // 1/148 = 0.0067567568
      10'd149: inv_x_count = 16'b0000000110111000; // 1/149 = 0.0067114094
      10'd150: inv_x_count = 16'b0000000110110101; // 1/150 = 0.0066666667
      10'd151: inv_x_count = 16'b0000000110110010; // 1/151 = 0.0066225166
      10'd152: inv_x_count = 16'b0000000110101111; // 1/152 = 0.0065789474
      10'd153: inv_x_count = 16'b0000000110101100; // 1/153 = 0.0065359477
      10'd154: inv_x_count = 16'b0000000110101010; // 1/154 = 0.0064935065
      10'd155: inv_x_count = 16'b0000000110100111; // 1/155 = 0.0064516129
      10'd156: inv_x_count = 16'b0000000110100100; // 1/156 = 0.0064102564
      10'd157: inv_x_count = 16'b0000000110100001; // 1/157 = 0.0063694268
      10'd158: inv_x_count = 16'b0000000110011111; // 1/158 = 0.0063291139
      10'd159: inv_x_count = 16'b0000000110011100; // 1/159 = 0.0062893082
      10'd160: inv_x_count = 16'b0000000110011010; // 1/160 = 0.0062500000
      10'd161: inv_x_count = 16'b0000000110010111; // 1/161 = 0.0062111801
      10'd162: inv_x_count = 16'b0000000110010101; // 1/162 = 0.0061728395
      10'd163: inv_x_count = 16'b0000000110010010; // 1/163 = 0.0061349693
      10'd164: inv_x_count = 16'b0000000110010000; // 1/164 = 0.0060975610
      10'd165: inv_x_count = 16'b0000000110001101; // 1/165 = 0.0060606061
      10'd166: inv_x_count = 16'b0000000110001011; // 1/166 = 0.0060240964
      10'd167: inv_x_count = 16'b0000000110001000; // 1/167 = 0.0059880240
      10'd168: inv_x_count = 16'b0000000110000110; // 1/168 = 0.0059523810
      10'd169: inv_x_count = 16'b0000000110000100; // 1/169 = 0.0059171598
      10'd170: inv_x_count = 16'b0000000110000010; // 1/170 = 0.0058823529
      10'd171: inv_x_count = 16'b0000000101111111; // 1/171 = 0.0058479532
      10'd172: inv_x_count = 16'b0000000101111101; // 1/172 = 0.0058139535
      10'd173: inv_x_count = 16'b0000000101111011; // 1/173 = 0.0057803468
      10'd174: inv_x_count = 16'b0000000101111001; // 1/174 = 0.0057471264
      10'd175: inv_x_count = 16'b0000000101110110; // 1/175 = 0.0057142857
      10'd176: inv_x_count = 16'b0000000101110100; // 1/176 = 0.0056818182
      10'd177: inv_x_count = 16'b0000000101110010; // 1/177 = 0.0056497175
      10'd178: inv_x_count = 16'b0000000101110000; // 1/178 = 0.0056179775
      10'd179: inv_x_count = 16'b0000000101101110; // 1/179 = 0.0055865922
      10'd180: inv_x_count = 16'b0000000101101100; // 1/180 = 0.0055555556
      10'd181: inv_x_count = 16'b0000000101101010; // 1/181 = 0.0055248619
      10'd182: inv_x_count = 16'b0000000101101000; // 1/182 = 0.0054945055
      10'd183: inv_x_count = 16'b0000000101100110; // 1/183 = 0.0054644809
      10'd184: inv_x_count = 16'b0000000101100100; // 1/184 = 0.0054347826
      10'd185: inv_x_count = 16'b0000000101100010; // 1/185 = 0.0054054054
      10'd186: inv_x_count = 16'b0000000101100000; // 1/186 = 0.0053763441
      10'd187: inv_x_count = 16'b0000000101011110; // 1/187 = 0.0053475936
      10'd188: inv_x_count = 16'b0000000101011101; // 1/188 = 0.0053191489
      10'd189: inv_x_count = 16'b0000000101011011; // 1/189 = 0.0052910053
      10'd190: inv_x_count = 16'b0000000101011001; // 1/190 = 0.0052631579
      10'd191: inv_x_count = 16'b0000000101010111; // 1/191 = 0.0052356021
      10'd192: inv_x_count = 16'b0000000101010101; // 1/192 = 0.0052083333
      10'd193: inv_x_count = 16'b0000000101010100; // 1/193 = 0.0051813472
      10'd194: inv_x_count = 16'b0000000101010010; // 1/194 = 0.0051546392
      10'd195: inv_x_count = 16'b0000000101010000; // 1/195 = 0.0051282051
      10'd196: inv_x_count = 16'b0000000101001110; // 1/196 = 0.0051020408
      10'd197: inv_x_count = 16'b0000000101001101; // 1/197 = 0.0050761421
      10'd198: inv_x_count = 16'b0000000101001011; // 1/198 = 0.0050505051
      10'd199: inv_x_count = 16'b0000000101001001; // 1/199 = 0.0050251256
      10'd200: inv_x_count = 16'b0000000101001000; // 1/200 = 0.0050000000
      10'd201: inv_x_count = 16'b0000000101000110; // 1/201 = 0.0049751244
      10'd202: inv_x_count = 16'b0000000101000100; // 1/202 = 0.0049504950
      10'd203: inv_x_count = 16'b0000000101000011; // 1/203 = 0.0049261084
      10'd204: inv_x_count = 16'b0000000101000001; // 1/204 = 0.0049019608
      10'd205: inv_x_count = 16'b0000000101000000; // 1/205 = 0.0048780488
      10'd206: inv_x_count = 16'b0000000100111110; // 1/206 = 0.0048543689
      10'd207: inv_x_count = 16'b0000000100111101; // 1/207 = 0.0048309179
      10'd208: inv_x_count = 16'b0000000100111011; // 1/208 = 0.0048076923
      10'd209: inv_x_count = 16'b0000000100111010; // 1/209 = 0.0047846890
      10'd210: inv_x_count = 16'b0000000100111000; // 1/210 = 0.0047619048
      10'd211: inv_x_count = 16'b0000000100110111; // 1/211 = 0.0047393365
      10'd212: inv_x_count = 16'b0000000100110101; // 1/212 = 0.0047169811
      10'd213: inv_x_count = 16'b0000000100110100; // 1/213 = 0.0046948357
      10'd214: inv_x_count = 16'b0000000100110010; // 1/214 = 0.0046728972
      10'd215: inv_x_count = 16'b0000000100110001; // 1/215 = 0.0046511628
      10'd216: inv_x_count = 16'b0000000100101111; // 1/216 = 0.0046296296
      10'd217: inv_x_count = 16'b0000000100101110; // 1/217 = 0.0046082949
      10'd218: inv_x_count = 16'b0000000100101101; // 1/218 = 0.0045871560
      10'd219: inv_x_count = 16'b0000000100101011; // 1/219 = 0.0045662100
      10'd220: inv_x_count = 16'b0000000100101010; // 1/220 = 0.0045454545
      10'd221: inv_x_count = 16'b0000000100101001; // 1/221 = 0.0045248869
      10'd222: inv_x_count = 16'b0000000100100111; // 1/222 = 0.0045045045
      10'd223: inv_x_count = 16'b0000000100100110; // 1/223 = 0.0044843049
      10'd224: inv_x_count = 16'b0000000100100101; // 1/224 = 0.0044642857
      10'd225: inv_x_count = 16'b0000000100100011; // 1/225 = 0.0044444444
      10'd226: inv_x_count = 16'b0000000100100010; // 1/226 = 0.0044247788
      10'd227: inv_x_count = 16'b0000000100100001; // 1/227 = 0.0044052863
      10'd228: inv_x_count = 16'b0000000100011111; // 1/228 = 0.0043859649
      10'd229: inv_x_count = 16'b0000000100011110; // 1/229 = 0.0043668122
      10'd230: inv_x_count = 16'b0000000100011101; // 1/230 = 0.0043478261
      10'd231: inv_x_count = 16'b0000000100011100; // 1/231 = 0.0043290043
      10'd232: inv_x_count = 16'b0000000100011010; // 1/232 = 0.0043103448
      10'd233: inv_x_count = 16'b0000000100011001; // 1/233 = 0.0042918455
      10'd234: inv_x_count = 16'b0000000100011000; // 1/234 = 0.0042735043
      10'd235: inv_x_count = 16'b0000000100010111; // 1/235 = 0.0042553191
      10'd236: inv_x_count = 16'b0000000100010110; // 1/236 = 0.0042372881
      10'd237: inv_x_count = 16'b0000000100010101; // 1/237 = 0.0042194093
      10'd238: inv_x_count = 16'b0000000100010011; // 1/238 = 0.0042016807
      10'd239: inv_x_count = 16'b0000000100010010; // 1/239 = 0.0041841004
      10'd240: inv_x_count = 16'b0000000100010001; // 1/240 = 0.0041666667
      10'd241: inv_x_count = 16'b0000000100010000; // 1/241 = 0.0041493776
      10'd242: inv_x_count = 16'b0000000100001111; // 1/242 = 0.0041322314
      10'd243: inv_x_count = 16'b0000000100001110; // 1/243 = 0.0041152263
      10'd244: inv_x_count = 16'b0000000100001101; // 1/244 = 0.0040983607
      10'd245: inv_x_count = 16'b0000000100001011; // 1/245 = 0.0040816327
      10'd246: inv_x_count = 16'b0000000100001010; // 1/246 = 0.0040650407
      10'd247: inv_x_count = 16'b0000000100001001; // 1/247 = 0.0040485830
      10'd248: inv_x_count = 16'b0000000100001000; // 1/248 = 0.0040322581
      10'd249: inv_x_count = 16'b0000000100000111; // 1/249 = 0.0040160643
      10'd250: inv_x_count = 16'b0000000100000110; // 1/250 = 0.0040000000
      10'd251: inv_x_count = 16'b0000000100000101; // 1/251 = 0.0039840637
      10'd252: inv_x_count = 16'b0000000100000100; // 1/252 = 0.0039682540
      10'd253: inv_x_count = 16'b0000000100000011; // 1/253 = 0.0039525692
      10'd254: inv_x_count = 16'b0000000100000010; // 1/254 = 0.0039370079
      10'd255: inv_x_count = 16'b0000000100000001; // 1/255 = 0.0039215686
      10'd256: inv_x_count = 16'b0000000100000000; // 1/256 = 0.0039062500
      10'd257: inv_x_count = 16'b0000000011111111; // 1/257 = 0.0038910506
      10'd258: inv_x_count = 16'b0000000011111110; // 1/258 = 0.0038759690
      10'd259: inv_x_count = 16'b0000000011111101; // 1/259 = 0.0038610039
      10'd260: inv_x_count = 16'b0000000011111100; // 1/260 = 0.0038461538
      10'd261: inv_x_count = 16'b0000000011111011; // 1/261 = 0.0038314176
      10'd262: inv_x_count = 16'b0000000011111010; // 1/262 = 0.0038167939
      10'd263: inv_x_count = 16'b0000000011111001; // 1/263 = 0.0038022814
      10'd264: inv_x_count = 16'b0000000011111000; // 1/264 = 0.0037878788
      10'd265: inv_x_count = 16'b0000000011110111; // 1/265 = 0.0037735849
      10'd266: inv_x_count = 16'b0000000011110110; // 1/266 = 0.0037593985
      10'd267: inv_x_count = 16'b0000000011110101; // 1/267 = 0.0037453184
      10'd268: inv_x_count = 16'b0000000011110101; // 1/268 = 0.0037313433
      10'd269: inv_x_count = 16'b0000000011110100; // 1/269 = 0.0037174721
      10'd270: inv_x_count = 16'b0000000011110011; // 1/270 = 0.0037037037
      10'd271: inv_x_count = 16'b0000000011110010; // 1/271 = 0.0036900369
      10'd272: inv_x_count = 16'b0000000011110001; // 1/272 = 0.0036764706
      10'd273: inv_x_count = 16'b0000000011110000; // 1/273 = 0.0036630037
      10'd274: inv_x_count = 16'b0000000011101111; // 1/274 = 0.0036496350
      10'd275: inv_x_count = 16'b0000000011101110; // 1/275 = 0.0036363636
      10'd276: inv_x_count = 16'b0000000011101101; // 1/276 = 0.0036231884
      10'd277: inv_x_count = 16'b0000000011101101; // 1/277 = 0.0036101083
      10'd278: inv_x_count = 16'b0000000011101100; // 1/278 = 0.0035971223
      10'd279: inv_x_count = 16'b0000000011101011; // 1/279 = 0.0035842294
      10'd280: inv_x_count = 16'b0000000011101010; // 1/280 = 0.0035714286
      10'd281: inv_x_count = 16'b0000000011101001; // 1/281 = 0.0035587189
      10'd282: inv_x_count = 16'b0000000011101000; // 1/282 = 0.0035460993
      10'd283: inv_x_count = 16'b0000000011101000; // 1/283 = 0.0035335689
      10'd284: inv_x_count = 16'b0000000011100111; // 1/284 = 0.0035211268
      10'd285: inv_x_count = 16'b0000000011100110; // 1/285 = 0.0035087719
      10'd286: inv_x_count = 16'b0000000011100101; // 1/286 = 0.0034965035
      10'd287: inv_x_count = 16'b0000000011100100; // 1/287 = 0.0034843206
      10'd288: inv_x_count = 16'b0000000011100100; // 1/288 = 0.0034722222
      10'd289: inv_x_count = 16'b0000000011100011; // 1/289 = 0.0034602076
      10'd290: inv_x_count = 16'b0000000011100010; // 1/290 = 0.0034482759
      10'd291: inv_x_count = 16'b0000000011100001; // 1/291 = 0.0034364261
      10'd292: inv_x_count = 16'b0000000011100000; // 1/292 = 0.0034246575
      10'd293: inv_x_count = 16'b0000000011100000; // 1/293 = 0.0034129693
      10'd294: inv_x_count = 16'b0000000011011111; // 1/294 = 0.0034013605
      10'd295: inv_x_count = 16'b0000000011011110; // 1/295 = 0.0033898305
      10'd296: inv_x_count = 16'b0000000011011101; // 1/296 = 0.0033783784
      10'd297: inv_x_count = 16'b0000000011011101; // 1/297 = 0.0033670034
      10'd298: inv_x_count = 16'b0000000011011100; // 1/298 = 0.0033557047
      10'd299: inv_x_count = 16'b0000000011011011; // 1/299 = 0.0033444816
      10'd300: inv_x_count = 16'b0000000011011010; // 1/300 = 0.0033333333
      10'd301: inv_x_count = 16'b0000000011011010; // 1/301 = 0.0033222591
      10'd302: inv_x_count = 16'b0000000011011001; // 1/302 = 0.0033112583
      10'd303: inv_x_count = 16'b0000000011011000; // 1/303 = 0.0033003300
      10'd304: inv_x_count = 16'b0000000011011000; // 1/304 = 0.0032894737
      10'd305: inv_x_count = 16'b0000000011010111; // 1/305 = 0.0032786885
      10'd306: inv_x_count = 16'b0000000011010110; // 1/306 = 0.0032679739
      10'd307: inv_x_count = 16'b0000000011010101; // 1/307 = 0.0032573290
      10'd308: inv_x_count = 16'b0000000011010101; // 1/308 = 0.0032467532
      10'd309: inv_x_count = 16'b0000000011010100; // 1/309 = 0.0032362460
      10'd310: inv_x_count = 16'b0000000011010011; // 1/310 = 0.0032258065
      10'd311: inv_x_count = 16'b0000000011010011; // 1/311 = 0.0032154341
      10'd312: inv_x_count = 16'b0000000011010010; // 1/312 = 0.0032051282
      10'd313: inv_x_count = 16'b0000000011010001; // 1/313 = 0.0031948882
      10'd314: inv_x_count = 16'b0000000011010001; // 1/314 = 0.0031847134
      10'd315: inv_x_count = 16'b0000000011010000; // 1/315 = 0.0031746032
      10'd316: inv_x_count = 16'b0000000011001111; // 1/316 = 0.0031645570
      10'd317: inv_x_count = 16'b0000000011001111; // 1/317 = 0.0031545741
      10'd318: inv_x_count = 16'b0000000011001110; // 1/318 = 0.0031446541
      10'd319: inv_x_count = 16'b0000000011001101; // 1/319 = 0.0031347962
      10'd320: inv_x_count = 16'b0000000011001101; // 1/320 = 0.0031250000
      10'd321: inv_x_count = 16'b0000000011001100; // 1/321 = 0.0031152648
      10'd322: inv_x_count = 16'b0000000011001100; // 1/322 = 0.0031055901
      10'd323: inv_x_count = 16'b0000000011001011; // 1/323 = 0.0030959752
      10'd324: inv_x_count = 16'b0000000011001010; // 1/324 = 0.0030864198
      10'd325: inv_x_count = 16'b0000000011001010; // 1/325 = 0.0030769231
      10'd326: inv_x_count = 16'b0000000011001001; // 1/326 = 0.0030674847
      10'd327: inv_x_count = 16'b0000000011001000; // 1/327 = 0.0030581040
      10'd328: inv_x_count = 16'b0000000011001000; // 1/328 = 0.0030487805
      10'd329: inv_x_count = 16'b0000000011000111; // 1/329 = 0.0030395137
      10'd330: inv_x_count = 16'b0000000011000111; // 1/330 = 0.0030303030
      10'd331: inv_x_count = 16'b0000000011000110; // 1/331 = 0.0030211480
      10'd332: inv_x_count = 16'b0000000011000101; // 1/332 = 0.0030120482
      10'd333: inv_x_count = 16'b0000000011000101; // 1/333 = 0.0030030030
      10'd334: inv_x_count = 16'b0000000011000100; // 1/334 = 0.0029940120
      10'd335: inv_x_count = 16'b0000000011000100; // 1/335 = 0.0029850746
      10'd336: inv_x_count = 16'b0000000011000011; // 1/336 = 0.0029761905
      10'd337: inv_x_count = 16'b0000000011000010; // 1/337 = 0.0029673591
      10'd338: inv_x_count = 16'b0000000011000010; // 1/338 = 0.0029585799
      10'd339: inv_x_count = 16'b0000000011000001; // 1/339 = 0.0029498525
      10'd340: inv_x_count = 16'b0000000011000001; // 1/340 = 0.0029411765
      10'd341: inv_x_count = 16'b0000000011000000; // 1/341 = 0.0029325513
      10'd342: inv_x_count = 16'b0000000011000000; // 1/342 = 0.0029239766
      10'd343: inv_x_count = 16'b0000000010111111; // 1/343 = 0.0029154519
      10'd344: inv_x_count = 16'b0000000010111111; // 1/344 = 0.0029069767
      10'd345: inv_x_count = 16'b0000000010111110; // 1/345 = 0.0028985507
      10'd346: inv_x_count = 16'b0000000010111101; // 1/346 = 0.0028901734
      10'd347: inv_x_count = 16'b0000000010111101; // 1/347 = 0.0028818444
      10'd348: inv_x_count = 16'b0000000010111100; // 1/348 = 0.0028735632
      10'd349: inv_x_count = 16'b0000000010111100; // 1/349 = 0.0028653295
      10'd350: inv_x_count = 16'b0000000010111011; // 1/350 = 0.0028571429
      10'd351: inv_x_count = 16'b0000000010111011; // 1/351 = 0.0028490028
      10'd352: inv_x_count = 16'b0000000010111010; // 1/352 = 0.0028409091
      10'd353: inv_x_count = 16'b0000000010111010; // 1/353 = 0.0028328612
      10'd354: inv_x_count = 16'b0000000010111001; // 1/354 = 0.0028248588
      10'd355: inv_x_count = 16'b0000000010111001; // 1/355 = 0.0028169014
      10'd356: inv_x_count = 16'b0000000010111000; // 1/356 = 0.0028089888
      10'd357: inv_x_count = 16'b0000000010111000; // 1/357 = 0.0028011204
      10'd358: inv_x_count = 16'b0000000010110111; // 1/358 = 0.0027932961
      10'd359: inv_x_count = 16'b0000000010110111; // 1/359 = 0.0027855153
      10'd360: inv_x_count = 16'b0000000010110110; // 1/360 = 0.0027777778
      10'd361: inv_x_count = 16'b0000000010110110; // 1/361 = 0.0027700831
      10'd362: inv_x_count = 16'b0000000010110101; // 1/362 = 0.0027624309
      10'd363: inv_x_count = 16'b0000000010110101; // 1/363 = 0.0027548209
      10'd364: inv_x_count = 16'b0000000010110100; // 1/364 = 0.0027472527
      10'd365: inv_x_count = 16'b0000000010110100; // 1/365 = 0.0027397260
      10'd366: inv_x_count = 16'b0000000010110011; // 1/366 = 0.0027322404
      10'd367: inv_x_count = 16'b0000000010110011; // 1/367 = 0.0027247956
      10'd368: inv_x_count = 16'b0000000010110010; // 1/368 = 0.0027173913
      10'd369: inv_x_count = 16'b0000000010110010; // 1/369 = 0.0027100271
      10'd370: inv_x_count = 16'b0000000010110001; // 1/370 = 0.0027027027
      10'd371: inv_x_count = 16'b0000000010110001; // 1/371 = 0.0026954178
      10'd372: inv_x_count = 16'b0000000010110000; // 1/372 = 0.0026881720
      10'd373: inv_x_count = 16'b0000000010110000; // 1/373 = 0.0026809651
      10'd374: inv_x_count = 16'b0000000010101111; // 1/374 = 0.0026737968
      10'd375: inv_x_count = 16'b0000000010101111; // 1/375 = 0.0026666667
      10'd376: inv_x_count = 16'b0000000010101110; // 1/376 = 0.0026595745
      10'd377: inv_x_count = 16'b0000000010101110; // 1/377 = 0.0026525199
      10'd378: inv_x_count = 16'b0000000010101101; // 1/378 = 0.0026455026
      10'd379: inv_x_count = 16'b0000000010101101; // 1/379 = 0.0026385224
      10'd380: inv_x_count = 16'b0000000010101100; // 1/380 = 0.0026315789
      10'd381: inv_x_count = 16'b0000000010101100; // 1/381 = 0.0026246719
      10'd382: inv_x_count = 16'b0000000010101100; // 1/382 = 0.0026178010
      10'd383: inv_x_count = 16'b0000000010101011; // 1/383 = 0.0026109661
      10'd384: inv_x_count = 16'b0000000010101011; // 1/384 = 0.0026041667
      10'd385: inv_x_count = 16'b0000000010101010; // 1/385 = 0.0025974026
      10'd386: inv_x_count = 16'b0000000010101010; // 1/386 = 0.0025906736
      10'd387: inv_x_count = 16'b0000000010101001; // 1/387 = 0.0025839793
      10'd388: inv_x_count = 16'b0000000010101001; // 1/388 = 0.0025773196
      10'd389: inv_x_count = 16'b0000000010101000; // 1/389 = 0.0025706941
      10'd390: inv_x_count = 16'b0000000010101000; // 1/390 = 0.0025641026
      10'd391: inv_x_count = 16'b0000000010101000; // 1/391 = 0.0025575448
      10'd392: inv_x_count = 16'b0000000010100111; // 1/392 = 0.0025510204
      10'd393: inv_x_count = 16'b0000000010100111; // 1/393 = 0.0025445293
      10'd394: inv_x_count = 16'b0000000010100110; // 1/394 = 0.0025380711
      10'd395: inv_x_count = 16'b0000000010100110; // 1/395 = 0.0025316456
      10'd396: inv_x_count = 16'b0000000010100101; // 1/396 = 0.0025252525
      10'd397: inv_x_count = 16'b0000000010100101; // 1/397 = 0.0025188917
      10'd398: inv_x_count = 16'b0000000010100101; // 1/398 = 0.0025125628
      10'd399: inv_x_count = 16'b0000000010100100; // 1/399 = 0.0025062657
      10'd400: inv_x_count = 16'b0000000010100100; // 1/400 = 0.0025000000
      10'd401: inv_x_count = 16'b0000000010100011; // 1/401 = 0.0024937656
      10'd402: inv_x_count = 16'b0000000010100011; // 1/402 = 0.0024875622
      10'd403: inv_x_count = 16'b0000000010100011; // 1/403 = 0.0024813896
      10'd404: inv_x_count = 16'b0000000010100010; // 1/404 = 0.0024752475
      10'd405: inv_x_count = 16'b0000000010100010; // 1/405 = 0.0024691358
      10'd406: inv_x_count = 16'b0000000010100001; // 1/406 = 0.0024630542
      10'd407: inv_x_count = 16'b0000000010100001; // 1/407 = 0.0024570025
      10'd408: inv_x_count = 16'b0000000010100001; // 1/408 = 0.0024509804
      10'd409: inv_x_count = 16'b0000000010100000; // 1/409 = 0.0024449878
      10'd410: inv_x_count = 16'b0000000010100000; // 1/410 = 0.0024390244
      10'd411: inv_x_count = 16'b0000000010011111; // 1/411 = 0.0024330900
      10'd412: inv_x_count = 16'b0000000010011111; // 1/412 = 0.0024271845
      10'd413: inv_x_count = 16'b0000000010011111; // 1/413 = 0.0024213075
      10'd414: inv_x_count = 16'b0000000010011110; // 1/414 = 0.0024154589
      10'd415: inv_x_count = 16'b0000000010011110; // 1/415 = 0.0024096386
      10'd416: inv_x_count = 16'b0000000010011110; // 1/416 = 0.0024038462
      10'd417: inv_x_count = 16'b0000000010011101; // 1/417 = 0.0023980815
      10'd418: inv_x_count = 16'b0000000010011101; // 1/418 = 0.0023923445
      10'd419: inv_x_count = 16'b0000000010011100; // 1/419 = 0.0023866348
      10'd420: inv_x_count = 16'b0000000010011100; // 1/420 = 0.0023809524
      10'd421: inv_x_count = 16'b0000000010011100; // 1/421 = 0.0023752969
      10'd422: inv_x_count = 16'b0000000010011011; // 1/422 = 0.0023696682
      10'd423: inv_x_count = 16'b0000000010011011; // 1/423 = 0.0023640662
      10'd424: inv_x_count = 16'b0000000010011011; // 1/424 = 0.0023584906
      10'd425: inv_x_count = 16'b0000000010011010; // 1/425 = 0.0023529412
      10'd426: inv_x_count = 16'b0000000010011010; // 1/426 = 0.0023474178
      10'd427: inv_x_count = 16'b0000000010011001; // 1/427 = 0.0023419204
      10'd428: inv_x_count = 16'b0000000010011001; // 1/428 = 0.0023364486
      10'd429: inv_x_count = 16'b0000000010011001; // 1/429 = 0.0023310023
      10'd430: inv_x_count = 16'b0000000010011000; // 1/430 = 0.0023255814
      10'd431: inv_x_count = 16'b0000000010011000; // 1/431 = 0.0023201856
      10'd432: inv_x_count = 16'b0000000010011000; // 1/432 = 0.0023148148
      10'd433: inv_x_count = 16'b0000000010010111; // 1/433 = 0.0023094688
      10'd434: inv_x_count = 16'b0000000010010111; // 1/434 = 0.0023041475
      10'd435: inv_x_count = 16'b0000000010010111; // 1/435 = 0.0022988506
      10'd436: inv_x_count = 16'b0000000010010110; // 1/436 = 0.0022935780
      10'd437: inv_x_count = 16'b0000000010010110; // 1/437 = 0.0022883295
      10'd438: inv_x_count = 16'b0000000010010110; // 1/438 = 0.0022831050
      10'd439: inv_x_count = 16'b0000000010010101; // 1/439 = 0.0022779043
      10'd440: inv_x_count = 16'b0000000010010101; // 1/440 = 0.0022727273
      10'd441: inv_x_count = 16'b0000000010010101; // 1/441 = 0.0022675737
      10'd442: inv_x_count = 16'b0000000010010100; // 1/442 = 0.0022624434
      10'd443: inv_x_count = 16'b0000000010010100; // 1/443 = 0.0022573363
      10'd444: inv_x_count = 16'b0000000010010100; // 1/444 = 0.0022522523
      10'd445: inv_x_count = 16'b0000000010010011; // 1/445 = 0.0022471910
      10'd446: inv_x_count = 16'b0000000010010011; // 1/446 = 0.0022421525
      10'd447: inv_x_count = 16'b0000000010010011; // 1/447 = 0.0022371365
      10'd448: inv_x_count = 16'b0000000010010010; // 1/448 = 0.0022321429
      10'd449: inv_x_count = 16'b0000000010010010; // 1/449 = 0.0022271715
      10'd450: inv_x_count = 16'b0000000010010010; // 1/450 = 0.0022222222
      10'd451: inv_x_count = 16'b0000000010010001; // 1/451 = 0.0022172949
      10'd452: inv_x_count = 16'b0000000010010001; // 1/452 = 0.0022123894
      10'd453: inv_x_count = 16'b0000000010010001; // 1/453 = 0.0022075055
      10'd454: inv_x_count = 16'b0000000010010000; // 1/454 = 0.0022026432
      10'd455: inv_x_count = 16'b0000000010010000; // 1/455 = 0.0021978022
      10'd456: inv_x_count = 16'b0000000010010000; // 1/456 = 0.0021929825
      10'd457: inv_x_count = 16'b0000000010001111; // 1/457 = 0.0021881838
      10'd458: inv_x_count = 16'b0000000010001111; // 1/458 = 0.0021834061
      10'd459: inv_x_count = 16'b0000000010001111; // 1/459 = 0.0021786492
      10'd460: inv_x_count = 16'b0000000010001110; // 1/460 = 0.0021739130
      10'd461: inv_x_count = 16'b0000000010001110; // 1/461 = 0.0021691974
      10'd462: inv_x_count = 16'b0000000010001110; // 1/462 = 0.0021645022
      10'd463: inv_x_count = 16'b0000000010001110; // 1/463 = 0.0021598272
      10'd464: inv_x_count = 16'b0000000010001101; // 1/464 = 0.0021551724
      10'd465: inv_x_count = 16'b0000000010001101; // 1/465 = 0.0021505376
      10'd466: inv_x_count = 16'b0000000010001101; // 1/466 = 0.0021459227
      10'd467: inv_x_count = 16'b0000000010001100; // 1/467 = 0.0021413276
      10'd468: inv_x_count = 16'b0000000010001100; // 1/468 = 0.0021367521
      10'd469: inv_x_count = 16'b0000000010001100; // 1/469 = 0.0021321962
      10'd470: inv_x_count = 16'b0000000010001011; // 1/470 = 0.0021276596
      10'd471: inv_x_count = 16'b0000000010001011; // 1/471 = 0.0021231423
      10'd472: inv_x_count = 16'b0000000010001011; // 1/472 = 0.0021186441
      10'd473: inv_x_count = 16'b0000000010001011; // 1/473 = 0.0021141649
      10'd474: inv_x_count = 16'b0000000010001010; // 1/474 = 0.0021097046
      10'd475: inv_x_count = 16'b0000000010001010; // 1/475 = 0.0021052632
      10'd476: inv_x_count = 16'b0000000010001010; // 1/476 = 0.0021008403
      10'd477: inv_x_count = 16'b0000000010001001; // 1/477 = 0.0020964361
      10'd478: inv_x_count = 16'b0000000010001001; // 1/478 = 0.0020920502
      10'd479: inv_x_count = 16'b0000000010001001; // 1/479 = 0.0020876827
      10'd480: inv_x_count = 16'b0000000010001001; // 1/480 = 0.0020833333
      10'd481: inv_x_count = 16'b0000000010001000; // 1/481 = 0.0020790021
      10'd482: inv_x_count = 16'b0000000010001000; // 1/482 = 0.0020746888
      10'd483: inv_x_count = 16'b0000000010001000; // 1/483 = 0.0020703934
      10'd484: inv_x_count = 16'b0000000010000111; // 1/484 = 0.0020661157
      10'd485: inv_x_count = 16'b0000000010000111; // 1/485 = 0.0020618557
      10'd486: inv_x_count = 16'b0000000010000111; // 1/486 = 0.0020576132
      10'd487: inv_x_count = 16'b0000000010000111; // 1/487 = 0.0020533881
      10'd488: inv_x_count = 16'b0000000010000110; // 1/488 = 0.0020491803
      10'd489: inv_x_count = 16'b0000000010000110; // 1/489 = 0.0020449898
      10'd490: inv_x_count = 16'b0000000010000110; // 1/490 = 0.0020408163
      10'd491: inv_x_count = 16'b0000000010000101; // 1/491 = 0.0020366599
      10'd492: inv_x_count = 16'b0000000010000101; // 1/492 = 0.0020325203
      10'd493: inv_x_count = 16'b0000000010000101; // 1/493 = 0.0020283976
      10'd494: inv_x_count = 16'b0000000010000101; // 1/494 = 0.0020242915
      10'd495: inv_x_count = 16'b0000000010000100; // 1/495 = 0.0020202020
      10'd496: inv_x_count = 16'b0000000010000100; // 1/496 = 0.0020161290
      10'd497: inv_x_count = 16'b0000000010000100; // 1/497 = 0.0020120724
      10'd498: inv_x_count = 16'b0000000010000100; // 1/498 = 0.0020080321
      10'd499: inv_x_count = 16'b0000000010000011; // 1/499 = 0.0020040080
      10'd500: inv_x_count = 16'b0000000010000011; // 1/500 = 0.0020000000
      10'd501: inv_x_count = 16'b0000000010000011; // 1/501 = 0.0019960080
      10'd502: inv_x_count = 16'b0000000010000011; // 1/502 = 0.0019920319
      10'd503: inv_x_count = 16'b0000000010000010; // 1/503 = 0.0019880716
      10'd504: inv_x_count = 16'b0000000010000010; // 1/504 = 0.0019841270
      10'd505: inv_x_count = 16'b0000000010000010; // 1/505 = 0.0019801980
      10'd506: inv_x_count = 16'b0000000010000010; // 1/506 = 0.0019762846
      10'd507: inv_x_count = 16'b0000000010000001; // 1/507 = 0.0019723866
      10'd508: inv_x_count = 16'b0000000010000001; // 1/508 = 0.0019685039
      10'd509: inv_x_count = 16'b0000000010000001; // 1/509 = 0.0019646365
      10'd510: inv_x_count = 16'b0000000010000001; // 1/510 = 0.0019607843
      10'd511: inv_x_count = 16'b0000000010000000; // 1/511 = 0.0019569472
      10'd512: inv_x_count = 16'b0000000010000000; // 1/512 = 0.0019531250
      10'd513: inv_x_count = 16'b0000000010000000; // 1/513 = 0.0019493177
      10'd514: inv_x_count = 16'b0000000010000000; // 1/514 = 0.0019455253
      10'd515: inv_x_count = 16'b0000000001111111; // 1/515 = 0.0019417476
      10'd516: inv_x_count = 16'b0000000001111111; // 1/516 = 0.0019379845
      10'd517: inv_x_count = 16'b0000000001111111; // 1/517 = 0.0019342360
      10'd518: inv_x_count = 16'b0000000001111111; // 1/518 = 0.0019305019
      10'd519: inv_x_count = 16'b0000000001111110; // 1/519 = 0.0019267823
      10'd520: inv_x_count = 16'b0000000001111110; // 1/520 = 0.0019230769
      10'd521: inv_x_count = 16'b0000000001111110; // 1/521 = 0.0019193858
      10'd522: inv_x_count = 16'b0000000001111110; // 1/522 = 0.0019157088
      10'd523: inv_x_count = 16'b0000000001111101; // 1/523 = 0.0019120459
      10'd524: inv_x_count = 16'b0000000001111101; // 1/524 = 0.0019083969
      10'd525: inv_x_count = 16'b0000000001111101; // 1/525 = 0.0019047619
      10'd526: inv_x_count = 16'b0000000001111101; // 1/526 = 0.0019011407
      10'd527: inv_x_count = 16'b0000000001111100; // 1/527 = 0.0018975332
      10'd528: inv_x_count = 16'b0000000001111100; // 1/528 = 0.0018939394
      10'd529: inv_x_count = 16'b0000000001111100; // 1/529 = 0.0018903592
      10'd530: inv_x_count = 16'b0000000001111100; // 1/530 = 0.0018867925
      10'd531: inv_x_count = 16'b0000000001111011; // 1/531 = 0.0018832392
      10'd532: inv_x_count = 16'b0000000001111011; // 1/532 = 0.0018796992
      10'd533: inv_x_count = 16'b0000000001111011; // 1/533 = 0.0018761726
      10'd534: inv_x_count = 16'b0000000001111011; // 1/534 = 0.0018726592
      10'd535: inv_x_count = 16'b0000000001111010; // 1/535 = 0.0018691589
      10'd536: inv_x_count = 16'b0000000001111010; // 1/536 = 0.0018656716
      10'd537: inv_x_count = 16'b0000000001111010; // 1/537 = 0.0018621974
      10'd538: inv_x_count = 16'b0000000001111010; // 1/538 = 0.0018587361
      10'd539: inv_x_count = 16'b0000000001111010; // 1/539 = 0.0018552876
      10'd540: inv_x_count = 16'b0000000001111001; // 1/540 = 0.0018518519
      10'd541: inv_x_count = 16'b0000000001111001; // 1/541 = 0.0018484288
      10'd542: inv_x_count = 16'b0000000001111001; // 1/542 = 0.0018450185
      10'd543: inv_x_count = 16'b0000000001111001; // 1/543 = 0.0018416206
      10'd544: inv_x_count = 16'b0000000001111000; // 1/544 = 0.0018382353
      10'd545: inv_x_count = 16'b0000000001111000; // 1/545 = 0.0018348624
      10'd546: inv_x_count = 16'b0000000001111000; // 1/546 = 0.0018315018
      10'd547: inv_x_count = 16'b0000000001111000; // 1/547 = 0.0018281536
      10'd548: inv_x_count = 16'b0000000001111000; // 1/548 = 0.0018248175
      10'd549: inv_x_count = 16'b0000000001110111; // 1/549 = 0.0018214936
      10'd550: inv_x_count = 16'b0000000001110111; // 1/550 = 0.0018181818
      10'd551: inv_x_count = 16'b0000000001110111; // 1/551 = 0.0018148820
      10'd552: inv_x_count = 16'b0000000001110111; // 1/552 = 0.0018115942
      10'd553: inv_x_count = 16'b0000000001110111; // 1/553 = 0.0018083183
      10'd554: inv_x_count = 16'b0000000001110110; // 1/554 = 0.0018050542
      10'd555: inv_x_count = 16'b0000000001110110; // 1/555 = 0.0018018018
      10'd556: inv_x_count = 16'b0000000001110110; // 1/556 = 0.0017985612
      10'd557: inv_x_count = 16'b0000000001110110; // 1/557 = 0.0017953321
      10'd558: inv_x_count = 16'b0000000001110101; // 1/558 = 0.0017921147
      10'd559: inv_x_count = 16'b0000000001110101; // 1/559 = 0.0017889088
      10'd560: inv_x_count = 16'b0000000001110101; // 1/560 = 0.0017857143
      10'd561: inv_x_count = 16'b0000000001110101; // 1/561 = 0.0017825312
      10'd562: inv_x_count = 16'b0000000001110101; // 1/562 = 0.0017793594
      10'd563: inv_x_count = 16'b0000000001110100; // 1/563 = 0.0017761989
      10'd564: inv_x_count = 16'b0000000001110100; // 1/564 = 0.0017730496
      10'd565: inv_x_count = 16'b0000000001110100; // 1/565 = 0.0017699115
      10'd566: inv_x_count = 16'b0000000001110100; // 1/566 = 0.0017667845
      10'd567: inv_x_count = 16'b0000000001110100; // 1/567 = 0.0017636684
      10'd568: inv_x_count = 16'b0000000001110011; // 1/568 = 0.0017605634
      10'd569: inv_x_count = 16'b0000000001110011; // 1/569 = 0.0017574692
      10'd570: inv_x_count = 16'b0000000001110011; // 1/570 = 0.0017543860
      10'd571: inv_x_count = 16'b0000000001110011; // 1/571 = 0.0017513135
      10'd572: inv_x_count = 16'b0000000001110011; // 1/572 = 0.0017482517
      10'd573: inv_x_count = 16'b0000000001110010; // 1/573 = 0.0017452007
      10'd574: inv_x_count = 16'b0000000001110010; // 1/574 = 0.0017421603
      10'd575: inv_x_count = 16'b0000000001110010; // 1/575 = 0.0017391304
      10'd576: inv_x_count = 16'b0000000001110010; // 1/576 = 0.0017361111
      10'd577: inv_x_count = 16'b0000000001110010; // 1/577 = 0.0017331023
      10'd578: inv_x_count = 16'b0000000001110001; // 1/578 = 0.0017301038
      10'd579: inv_x_count = 16'b0000000001110001; // 1/579 = 0.0017271157
      10'd580: inv_x_count = 16'b0000000001110001; // 1/580 = 0.0017241379
      10'd581: inv_x_count = 16'b0000000001110001; // 1/581 = 0.0017211704
      10'd582: inv_x_count = 16'b0000000001110001; // 1/582 = 0.0017182131
      10'd583: inv_x_count = 16'b0000000001110000; // 1/583 = 0.0017152659
      10'd584: inv_x_count = 16'b0000000001110000; // 1/584 = 0.0017123288
      10'd585: inv_x_count = 16'b0000000001110000; // 1/585 = 0.0017094017
      10'd586: inv_x_count = 16'b0000000001110000; // 1/586 = 0.0017064846
      10'd587: inv_x_count = 16'b0000000001110000; // 1/587 = 0.0017035775
      10'd588: inv_x_count = 16'b0000000001101111; // 1/588 = 0.0017006803
      10'd589: inv_x_count = 16'b0000000001101111; // 1/589 = 0.0016977929
      10'd590: inv_x_count = 16'b0000000001101111; // 1/590 = 0.0016949153
      10'd591: inv_x_count = 16'b0000000001101111; // 1/591 = 0.0016920474
      10'd592: inv_x_count = 16'b0000000001101111; // 1/592 = 0.0016891892
      10'd593: inv_x_count = 16'b0000000001101111; // 1/593 = 0.0016863406
      10'd594: inv_x_count = 16'b0000000001101110; // 1/594 = 0.0016835017
      10'd595: inv_x_count = 16'b0000000001101110; // 1/595 = 0.0016806723
      10'd596: inv_x_count = 16'b0000000001101110; // 1/596 = 0.0016778523
      10'd597: inv_x_count = 16'b0000000001101110; // 1/597 = 0.0016750419
      10'd598: inv_x_count = 16'b0000000001101110; // 1/598 = 0.0016722408
      10'd599: inv_x_count = 16'b0000000001101101; // 1/599 = 0.0016694491
      10'd600: inv_x_count = 16'b0000000001101101; // 1/600 = 0.0016666667
      10'd601: inv_x_count = 16'b0000000001101101; // 1/601 = 0.0016638935
      10'd602: inv_x_count = 16'b0000000001101101; // 1/602 = 0.0016611296
      10'd603: inv_x_count = 16'b0000000001101101; // 1/603 = 0.0016583748
      10'd604: inv_x_count = 16'b0000000001101101; // 1/604 = 0.0016556291
      10'd605: inv_x_count = 16'b0000000001101100; // 1/605 = 0.0016528926
      10'd606: inv_x_count = 16'b0000000001101100; // 1/606 = 0.0016501650
      10'd607: inv_x_count = 16'b0000000001101100; // 1/607 = 0.0016474465
      10'd608: inv_x_count = 16'b0000000001101100; // 1/608 = 0.0016447368
      10'd609: inv_x_count = 16'b0000000001101100; // 1/609 = 0.0016420361
      10'd610: inv_x_count = 16'b0000000001101011; // 1/610 = 0.0016393443
      10'd611: inv_x_count = 16'b0000000001101011; // 1/611 = 0.0016366612
      10'd612: inv_x_count = 16'b0000000001101011; // 1/612 = 0.0016339869
      10'd613: inv_x_count = 16'b0000000001101011; // 1/613 = 0.0016313214
      10'd614: inv_x_count = 16'b0000000001101011; // 1/614 = 0.0016286645
      10'd615: inv_x_count = 16'b0000000001101011; // 1/615 = 0.0016260163
      10'd616: inv_x_count = 16'b0000000001101010; // 1/616 = 0.0016233766
      10'd617: inv_x_count = 16'b0000000001101010; // 1/617 = 0.0016207455
      10'd618: inv_x_count = 16'b0000000001101010; // 1/618 = 0.0016181230
      10'd619: inv_x_count = 16'b0000000001101010; // 1/619 = 0.0016155089
      10'd620: inv_x_count = 16'b0000000001101010; // 1/620 = 0.0016129032
      10'd621: inv_x_count = 16'b0000000001101010; // 1/621 = 0.0016103060
      10'd622: inv_x_count = 16'b0000000001101001; // 1/622 = 0.0016077170
      10'd623: inv_x_count = 16'b0000000001101001; // 1/623 = 0.0016051364
      10'd624: inv_x_count = 16'b0000000001101001; // 1/624 = 0.0016025641
      10'd625: inv_x_count = 16'b0000000001101001; // 1/625 = 0.0016000000
      10'd626: inv_x_count = 16'b0000000001101001; // 1/626 = 0.0015974441
      10'd627: inv_x_count = 16'b0000000001101001; // 1/627 = 0.0015948963
      10'd628: inv_x_count = 16'b0000000001101000; // 1/628 = 0.0015923567
      10'd629: inv_x_count = 16'b0000000001101000; // 1/629 = 0.0015898251
      10'd630: inv_x_count = 16'b0000000001101000; // 1/630 = 0.0015873016
      10'd631: inv_x_count = 16'b0000000001101000; // 1/631 = 0.0015847861
      10'd632: inv_x_count = 16'b0000000001101000; // 1/632 = 0.0015822785
      10'd633: inv_x_count = 16'b0000000001101000; // 1/633 = 0.0015797788
      10'd634: inv_x_count = 16'b0000000001100111; // 1/634 = 0.0015772871
      10'd635: inv_x_count = 16'b0000000001100111; // 1/635 = 0.0015748031
      10'd636: inv_x_count = 16'b0000000001100111; // 1/636 = 0.0015723270
      10'd637: inv_x_count = 16'b0000000001100111; // 1/637 = 0.0015698587
      10'd638: inv_x_count = 16'b0000000001100111; // 1/638 = 0.0015673981
      10'd639: inv_x_count = 16'b0000000001100111; // 1/639 = 0.0015649452
      10'd640: inv_x_count = 16'b0000000001100110; // 1/640 = 0.0015625000
      10'd641: inv_x_count = 16'b0000000001100110; // 1/641 = 0.0015600624
      10'd642: inv_x_count = 16'b0000000001100110; // 1/642 = 0.0015576324
      10'd643: inv_x_count = 16'b0000000001100110; // 1/643 = 0.0015552100
      10'd644: inv_x_count = 16'b0000000001100110; // 1/644 = 0.0015527950
      10'd645: inv_x_count = 16'b0000000001100110; // 1/645 = 0.0015503876
      10'd646: inv_x_count = 16'b0000000001100101; // 1/646 = 0.0015479876
      10'd647: inv_x_count = 16'b0000000001100101; // 1/647 = 0.0015455951
      10'd648: inv_x_count = 16'b0000000001100101; // 1/648 = 0.0015432099
      10'd649: inv_x_count = 16'b0000000001100101; // 1/649 = 0.0015408320
      10'd650: inv_x_count = 16'b0000000001100101; // 1/650 = 0.0015384615
      10'd651: inv_x_count = 16'b0000000001100101; // 1/651 = 0.0015360983
      10'd652: inv_x_count = 16'b0000000001100101; // 1/652 = 0.0015337423
      10'd653: inv_x_count = 16'b0000000001100100; // 1/653 = 0.0015313936
      10'd654: inv_x_count = 16'b0000000001100100; // 1/654 = 0.0015290520
      10'd655: inv_x_count = 16'b0000000001100100; // 1/655 = 0.0015267176
      10'd656: inv_x_count = 16'b0000000001100100; // 1/656 = 0.0015243902
      10'd657: inv_x_count = 16'b0000000001100100; // 1/657 = 0.0015220700
      10'd658: inv_x_count = 16'b0000000001100100; // 1/658 = 0.0015197568
      10'd659: inv_x_count = 16'b0000000001100011; // 1/659 = 0.0015174507
      10'd660: inv_x_count = 16'b0000000001100011; // 1/660 = 0.0015151515
      10'd661: inv_x_count = 16'b0000000001100011; // 1/661 = 0.0015128593
      10'd662: inv_x_count = 16'b0000000001100011; // 1/662 = 0.0015105740
      10'd663: inv_x_count = 16'b0000000001100011; // 1/663 = 0.0015082956
      10'd664: inv_x_count = 16'b0000000001100011; // 1/664 = 0.0015060241
      10'd665: inv_x_count = 16'b0000000001100011; // 1/665 = 0.0015037594
      10'd666: inv_x_count = 16'b0000000001100010; // 1/666 = 0.0015015015
      10'd667: inv_x_count = 16'b0000000001100010; // 1/667 = 0.0014992504
      10'd668: inv_x_count = 16'b0000000001100010; // 1/668 = 0.0014970060
      10'd669: inv_x_count = 16'b0000000001100010; // 1/669 = 0.0014947683
      10'd670: inv_x_count = 16'b0000000001100010; // 1/670 = 0.0014925373
      10'd671: inv_x_count = 16'b0000000001100010; // 1/671 = 0.0014903130
      10'd672: inv_x_count = 16'b0000000001100010; // 1/672 = 0.0014880952
      10'd673: inv_x_count = 16'b0000000001100001; // 1/673 = 0.0014858841
      10'd674: inv_x_count = 16'b0000000001100001; // 1/674 = 0.0014836795
      10'd675: inv_x_count = 16'b0000000001100001; // 1/675 = 0.0014814815
      10'd676: inv_x_count = 16'b0000000001100001; // 1/676 = 0.0014792899
      10'd677: inv_x_count = 16'b0000000001100001; // 1/677 = 0.0014771049
      10'd678: inv_x_count = 16'b0000000001100001; // 1/678 = 0.0014749263
      10'd679: inv_x_count = 16'b0000000001100001; // 1/679 = 0.0014727541
      10'd680: inv_x_count = 16'b0000000001100000; // 1/680 = 0.0014705882
      10'd681: inv_x_count = 16'b0000000001100000; // 1/681 = 0.0014684288
      10'd682: inv_x_count = 16'b0000000001100000; // 1/682 = 0.0014662757
      10'd683: inv_x_count = 16'b0000000001100000; // 1/683 = 0.0014641288
      10'd684: inv_x_count = 16'b0000000001100000; // 1/684 = 0.0014619883
      10'd685: inv_x_count = 16'b0000000001100000; // 1/685 = 0.0014598540
      10'd686: inv_x_count = 16'b0000000001100000; // 1/686 = 0.0014577259
      10'd687: inv_x_count = 16'b0000000001011111; // 1/687 = 0.0014556041
      10'd688: inv_x_count = 16'b0000000001011111; // 1/688 = 0.0014534884
      10'd689: inv_x_count = 16'b0000000001011111; // 1/689 = 0.0014513788
      10'd690: inv_x_count = 16'b0000000001011111; // 1/690 = 0.0014492754
      10'd691: inv_x_count = 16'b0000000001011111; // 1/691 = 0.0014471780
      10'd692: inv_x_count = 16'b0000000001011111; // 1/692 = 0.0014450867
      10'd693: inv_x_count = 16'b0000000001011111; // 1/693 = 0.0014430014
      10'd694: inv_x_count = 16'b0000000001011110; // 1/694 = 0.0014409222
      10'd695: inv_x_count = 16'b0000000001011110; // 1/695 = 0.0014388489
      10'd696: inv_x_count = 16'b0000000001011110; // 1/696 = 0.0014367816
      10'd697: inv_x_count = 16'b0000000001011110; // 1/697 = 0.0014347202
      10'd698: inv_x_count = 16'b0000000001011110; // 1/698 = 0.0014326648
      10'd699: inv_x_count = 16'b0000000001011110; // 1/699 = 0.0014306152
      10'd700: inv_x_count = 16'b0000000001011110; // 1/700 = 0.0014285714
      10'd701: inv_x_count = 16'b0000000001011101; // 1/701 = 0.0014265335
      10'd702: inv_x_count = 16'b0000000001011101; // 1/702 = 0.0014245014
      10'd703: inv_x_count = 16'b0000000001011101; // 1/703 = 0.0014224751
      10'd704: inv_x_count = 16'b0000000001011101; // 1/704 = 0.0014204545
      10'd705: inv_x_count = 16'b0000000001011101; // 1/705 = 0.0014184397
      10'd706: inv_x_count = 16'b0000000001011101; // 1/706 = 0.0014164306
      10'd707: inv_x_count = 16'b0000000001011101; // 1/707 = 0.0014144272
      10'd708: inv_x_count = 16'b0000000001011101; // 1/708 = 0.0014124294
      10'd709: inv_x_count = 16'b0000000001011100; // 1/709 = 0.0014104372
      10'd710: inv_x_count = 16'b0000000001011100; // 1/710 = 0.0014084507
      10'd711: inv_x_count = 16'b0000000001011100; // 1/711 = 0.0014064698
      10'd712: inv_x_count = 16'b0000000001011100; // 1/712 = 0.0014044944
      10'd713: inv_x_count = 16'b0000000001011100; // 1/713 = 0.0014025245
      10'd714: inv_x_count = 16'b0000000001011100; // 1/714 = 0.0014005602
      10'd715: inv_x_count = 16'b0000000001011100; // 1/715 = 0.0013986014
      10'd716: inv_x_count = 16'b0000000001011100; // 1/716 = 0.0013966480
      10'd717: inv_x_count = 16'b0000000001011011; // 1/717 = 0.0013947001
      10'd718: inv_x_count = 16'b0000000001011011; // 1/718 = 0.0013927577
      10'd719: inv_x_count = 16'b0000000001011011; // 1/719 = 0.0013908206
      10'd720: inv_x_count = 16'b0000000001011011; // 1/720 = 0.0013888889
      10'd721: inv_x_count = 16'b0000000001011011; // 1/721 = 0.0013869626
      10'd722: inv_x_count = 16'b0000000001011011; // 1/722 = 0.0013850416
      10'd723: inv_x_count = 16'b0000000001011011; // 1/723 = 0.0013831259
      10'd724: inv_x_count = 16'b0000000001011011; // 1/724 = 0.0013812155
      10'd725: inv_x_count = 16'b0000000001011010; // 1/725 = 0.0013793103
      10'd726: inv_x_count = 16'b0000000001011010; // 1/726 = 0.0013774105
      10'd727: inv_x_count = 16'b0000000001011010; // 1/727 = 0.0013755158
      10'd728: inv_x_count = 16'b0000000001011010; // 1/728 = 0.0013736264
      10'd729: inv_x_count = 16'b0000000001011010; // 1/729 = 0.0013717421
      10'd730: inv_x_count = 16'b0000000001011010; // 1/730 = 0.0013698630
      10'd731: inv_x_count = 16'b0000000001011010; // 1/731 = 0.0013679891
      10'd732: inv_x_count = 16'b0000000001011010; // 1/732 = 0.0013661202
      10'd733: inv_x_count = 16'b0000000001011001; // 1/733 = 0.0013642565
      10'd734: inv_x_count = 16'b0000000001011001; // 1/734 = 0.0013623978
      10'd735: inv_x_count = 16'b0000000001011001; // 1/735 = 0.0013605442
      10'd736: inv_x_count = 16'b0000000001011001; // 1/736 = 0.0013586957
      10'd737: inv_x_count = 16'b0000000001011001; // 1/737 = 0.0013568521
      10'd738: inv_x_count = 16'b0000000001011001; // 1/738 = 0.0013550136
      10'd739: inv_x_count = 16'b0000000001011001; // 1/739 = 0.0013531800
      10'd740: inv_x_count = 16'b0000000001011001; // 1/740 = 0.0013513514
      10'd741: inv_x_count = 16'b0000000001011000; // 1/741 = 0.0013495277
      10'd742: inv_x_count = 16'b0000000001011000; // 1/742 = 0.0013477089
      10'd743: inv_x_count = 16'b0000000001011000; // 1/743 = 0.0013458950
      10'd744: inv_x_count = 16'b0000000001011000; // 1/744 = 0.0013440860
      10'd745: inv_x_count = 16'b0000000001011000; // 1/745 = 0.0013422819
      10'd746: inv_x_count = 16'b0000000001011000; // 1/746 = 0.0013404826
      10'd747: inv_x_count = 16'b0000000001011000; // 1/747 = 0.0013386881
      10'd748: inv_x_count = 16'b0000000001011000; // 1/748 = 0.0013368984
      10'd749: inv_x_count = 16'b0000000001010111; // 1/749 = 0.0013351135
      10'd750: inv_x_count = 16'b0000000001010111; // 1/750 = 0.0013333333
      10'd751: inv_x_count = 16'b0000000001010111; // 1/751 = 0.0013315579
      10'd752: inv_x_count = 16'b0000000001010111; // 1/752 = 0.0013297872
      10'd753: inv_x_count = 16'b0000000001010111; // 1/753 = 0.0013280212
      10'd754: inv_x_count = 16'b0000000001010111; // 1/754 = 0.0013262599
      10'd755: inv_x_count = 16'b0000000001010111; // 1/755 = 0.0013245033
      10'd756: inv_x_count = 16'b0000000001010111; // 1/756 = 0.0013227513
      10'd757: inv_x_count = 16'b0000000001010111; // 1/757 = 0.0013210040
      10'd758: inv_x_count = 16'b0000000001010110; // 1/758 = 0.0013192612
      10'd759: inv_x_count = 16'b0000000001010110; // 1/759 = 0.0013175231
      10'd760: inv_x_count = 16'b0000000001010110; // 1/760 = 0.0013157895
      10'd761: inv_x_count = 16'b0000000001010110; // 1/761 = 0.0013140604
      10'd762: inv_x_count = 16'b0000000001010110; // 1/762 = 0.0013123360
      10'd763: inv_x_count = 16'b0000000001010110; // 1/763 = 0.0013106160
      10'd764: inv_x_count = 16'b0000000001010110; // 1/764 = 0.0013089005
      10'd765: inv_x_count = 16'b0000000001010110; // 1/765 = 0.0013071895
      10'd766: inv_x_count = 16'b0000000001010110; // 1/766 = 0.0013054830
      10'd767: inv_x_count = 16'b0000000001010101; // 1/767 = 0.0013037810
      10'd768: inv_x_count = 16'b0000000001010101; // 1/768 = 0.0013020833
      10'd769: inv_x_count = 16'b0000000001010101; // 1/769 = 0.0013003901
      10'd770: inv_x_count = 16'b0000000001010101; // 1/770 = 0.0012987013
      10'd771: inv_x_count = 16'b0000000001010101; // 1/771 = 0.0012970169
      10'd772: inv_x_count = 16'b0000000001010101; // 1/772 = 0.0012953368
      10'd773: inv_x_count = 16'b0000000001010101; // 1/773 = 0.0012936611
      10'd774: inv_x_count = 16'b0000000001010101; // 1/774 = 0.0012919897
      10'd775: inv_x_count = 16'b0000000001010101; // 1/775 = 0.0012903226
      10'd776: inv_x_count = 16'b0000000001010100; // 1/776 = 0.0012886598
      10'd777: inv_x_count = 16'b0000000001010100; // 1/777 = 0.0012870013
      10'd778: inv_x_count = 16'b0000000001010100; // 1/778 = 0.0012853470
      10'd779: inv_x_count = 16'b0000000001010100; // 1/779 = 0.0012836970
      10'd780: inv_x_count = 16'b0000000001010100; // 1/780 = 0.0012820513
      10'd781: inv_x_count = 16'b0000000001010100; // 1/781 = 0.0012804097
      10'd782: inv_x_count = 16'b0000000001010100; // 1/782 = 0.0012787724
      10'd783: inv_x_count = 16'b0000000001010100; // 1/783 = 0.0012771392
      10'd784: inv_x_count = 16'b0000000001010100; // 1/784 = 0.0012755102
      10'd785: inv_x_count = 16'b0000000001010011; // 1/785 = 0.0012738854
      10'd786: inv_x_count = 16'b0000000001010011; // 1/786 = 0.0012722646
      10'd787: inv_x_count = 16'b0000000001010011; // 1/787 = 0.0012706480
      10'd788: inv_x_count = 16'b0000000001010011; // 1/788 = 0.0012690355
      10'd789: inv_x_count = 16'b0000000001010011; // 1/789 = 0.0012674271
      10'd790: inv_x_count = 16'b0000000001010011; // 1/790 = 0.0012658228
      10'd791: inv_x_count = 16'b0000000001010011; // 1/791 = 0.0012642225
      10'd792: inv_x_count = 16'b0000000001010011; // 1/792 = 0.0012626263
      10'd793: inv_x_count = 16'b0000000001010011; // 1/793 = 0.0012610340
      10'd794: inv_x_count = 16'b0000000001010011; // 1/794 = 0.0012594458
      10'd795: inv_x_count = 16'b0000000001010010; // 1/795 = 0.0012578616
      10'd796: inv_x_count = 16'b0000000001010010; // 1/796 = 0.0012562814
      10'd797: inv_x_count = 16'b0000000001010010; // 1/797 = 0.0012547051
      10'd798: inv_x_count = 16'b0000000001010010; // 1/798 = 0.0012531328
      10'd799: inv_x_count = 16'b0000000001010010; // 1/799 = 0.0012515645
      10'd800: inv_x_count = 16'b0000000001010010; // 1/800 = 0.0012500000
      10'd801: inv_x_count = 16'b0000000001010010; // 1/801 = 0.0012484395
      10'd802: inv_x_count = 16'b0000000001010010; // 1/802 = 0.0012468828
      10'd803: inv_x_count = 16'b0000000001010010; // 1/803 = 0.0012453300
      10'd804: inv_x_count = 16'b0000000001010010; // 1/804 = 0.0012437811
      10'd805: inv_x_count = 16'b0000000001010001; // 1/805 = 0.0012422360
      10'd806: inv_x_count = 16'b0000000001010001; // 1/806 = 0.0012406948
      10'd807: inv_x_count = 16'b0000000001010001; // 1/807 = 0.0012391574
      10'd808: inv_x_count = 16'b0000000001010001; // 1/808 = 0.0012376238
      10'd809: inv_x_count = 16'b0000000001010001; // 1/809 = 0.0012360939
      10'd810: inv_x_count = 16'b0000000001010001; // 1/810 = 0.0012345679
      10'd811: inv_x_count = 16'b0000000001010001; // 1/811 = 0.0012330456
      10'd812: inv_x_count = 16'b0000000001010001; // 1/812 = 0.0012315271
      10'd813: inv_x_count = 16'b0000000001010001; // 1/813 = 0.0012300123
      10'd814: inv_x_count = 16'b0000000001010001; // 1/814 = 0.0012285012
      10'd815: inv_x_count = 16'b0000000001010000; // 1/815 = 0.0012269939
      10'd816: inv_x_count = 16'b0000000001010000; // 1/816 = 0.0012254902
      10'd817: inv_x_count = 16'b0000000001010000; // 1/817 = 0.0012239902
      10'd818: inv_x_count = 16'b0000000001010000; // 1/818 = 0.0012224939
      10'd819: inv_x_count = 16'b0000000001010000; // 1/819 = 0.0012210012
      10'd820: inv_x_count = 16'b0000000001010000; // 1/820 = 0.0012195122
      10'd821: inv_x_count = 16'b0000000001010000; // 1/821 = 0.0012180268
      10'd822: inv_x_count = 16'b0000000001010000; // 1/822 = 0.0012165450
      10'd823: inv_x_count = 16'b0000000001010000; // 1/823 = 0.0012150668
      10'd824: inv_x_count = 16'b0000000001010000; // 1/824 = 0.0012135922
      10'd825: inv_x_count = 16'b0000000001001111; // 1/825 = 0.0012121212
      10'd826: inv_x_count = 16'b0000000001001111; // 1/826 = 0.0012106538
      10'd827: inv_x_count = 16'b0000000001001111; // 1/827 = 0.0012091898
      10'd828: inv_x_count = 16'b0000000001001111; // 1/828 = 0.0012077295
      10'd829: inv_x_count = 16'b0000000001001111; // 1/829 = 0.0012062726
      10'd830: inv_x_count = 16'b0000000001001111; // 1/830 = 0.0012048193
      10'd831: inv_x_count = 16'b0000000001001111; // 1/831 = 0.0012033694
      10'd832: inv_x_count = 16'b0000000001001111; // 1/832 = 0.0012019231
      10'd833: inv_x_count = 16'b0000000001001111; // 1/833 = 0.0012004802
      10'd834: inv_x_count = 16'b0000000001001111; // 1/834 = 0.0011990408
      10'd835: inv_x_count = 16'b0000000001001110; // 1/835 = 0.0011976048
      10'd836: inv_x_count = 16'b0000000001001110; // 1/836 = 0.0011961722
      10'd837: inv_x_count = 16'b0000000001001110; // 1/837 = 0.0011947431
      10'd838: inv_x_count = 16'b0000000001001110; // 1/838 = 0.0011933174
      10'd839: inv_x_count = 16'b0000000001001110; // 1/839 = 0.0011918951
      10'd840: inv_x_count = 16'b0000000001001110; // 1/840 = 0.0011904762
      10'd841: inv_x_count = 16'b0000000001001110; // 1/841 = 0.0011890606
      10'd842: inv_x_count = 16'b0000000001001110; // 1/842 = 0.0011876485
      10'd843: inv_x_count = 16'b0000000001001110; // 1/843 = 0.0011862396
      10'd844: inv_x_count = 16'b0000000001001110; // 1/844 = 0.0011848341
      10'd845: inv_x_count = 16'b0000000001001110; // 1/845 = 0.0011834320
      10'd846: inv_x_count = 16'b0000000001001101; // 1/846 = 0.0011820331
      10'd847: inv_x_count = 16'b0000000001001101; // 1/847 = 0.0011806375
      10'd848: inv_x_count = 16'b0000000001001101; // 1/848 = 0.0011792453
      10'd849: inv_x_count = 16'b0000000001001101; // 1/849 = 0.0011778563
      10'd850: inv_x_count = 16'b0000000001001101; // 1/850 = 0.0011764706
      10'd851: inv_x_count = 16'b0000000001001101; // 1/851 = 0.0011750881
      10'd852: inv_x_count = 16'b0000000001001101; // 1/852 = 0.0011737089
      10'd853: inv_x_count = 16'b0000000001001101; // 1/853 = 0.0011723329
      10'd854: inv_x_count = 16'b0000000001001101; // 1/854 = 0.0011709602
      10'd855: inv_x_count = 16'b0000000001001101; // 1/855 = 0.0011695906
      10'd856: inv_x_count = 16'b0000000001001101; // 1/856 = 0.0011682243
      10'd857: inv_x_count = 16'b0000000001001100; // 1/857 = 0.0011668611
      10'd858: inv_x_count = 16'b0000000001001100; // 1/858 = 0.0011655012
      10'd859: inv_x_count = 16'b0000000001001100; // 1/859 = 0.0011641444
      10'd860: inv_x_count = 16'b0000000001001100; // 1/860 = 0.0011627907
      10'd861: inv_x_count = 16'b0000000001001100; // 1/861 = 0.0011614402
      10'd862: inv_x_count = 16'b0000000001001100; // 1/862 = 0.0011600928
      10'd863: inv_x_count = 16'b0000000001001100; // 1/863 = 0.0011587486
      10'd864: inv_x_count = 16'b0000000001001100; // 1/864 = 0.0011574074
      10'd865: inv_x_count = 16'b0000000001001100; // 1/865 = 0.0011560694
      10'd866: inv_x_count = 16'b0000000001001100; // 1/866 = 0.0011547344
      10'd867: inv_x_count = 16'b0000000001001100; // 1/867 = 0.0011534025
      10'd868: inv_x_count = 16'b0000000001001100; // 1/868 = 0.0011520737
      10'd869: inv_x_count = 16'b0000000001001011; // 1/869 = 0.0011507480
      10'd870: inv_x_count = 16'b0000000001001011; // 1/870 = 0.0011494253
      10'd871: inv_x_count = 16'b0000000001001011; // 1/871 = 0.0011481056
      10'd872: inv_x_count = 16'b0000000001001011; // 1/872 = 0.0011467890
      10'd873: inv_x_count = 16'b0000000001001011; // 1/873 = 0.0011454754
      10'd874: inv_x_count = 16'b0000000001001011; // 1/874 = 0.0011441648
      10'd875: inv_x_count = 16'b0000000001001011; // 1/875 = 0.0011428571
      10'd876: inv_x_count = 16'b0000000001001011; // 1/876 = 0.0011415525
      10'd877: inv_x_count = 16'b0000000001001011; // 1/877 = 0.0011402509
      10'd878: inv_x_count = 16'b0000000001001011; // 1/878 = 0.0011389522
      10'd879: inv_x_count = 16'b0000000001001011; // 1/879 = 0.0011376564
      10'd880: inv_x_count = 16'b0000000001001010; // 1/880 = 0.0011363636
      10'd881: inv_x_count = 16'b0000000001001010; // 1/881 = 0.0011350738
      10'd882: inv_x_count = 16'b0000000001001010; // 1/882 = 0.0011337868
      10'd883: inv_x_count = 16'b0000000001001010; // 1/883 = 0.0011325028
      10'd884: inv_x_count = 16'b0000000001001010; // 1/884 = 0.0011312217
      10'd885: inv_x_count = 16'b0000000001001010; // 1/885 = 0.0011299435
      10'd886: inv_x_count = 16'b0000000001001010; // 1/886 = 0.0011286682
      10'd887: inv_x_count = 16'b0000000001001010; // 1/887 = 0.0011273957
      10'd888: inv_x_count = 16'b0000000001001010; // 1/888 = 0.0011261261
      10'd889: inv_x_count = 16'b0000000001001010; // 1/889 = 0.0011248594
      10'd890: inv_x_count = 16'b0000000001001010; // 1/890 = 0.0011235955
      10'd891: inv_x_count = 16'b0000000001001010; // 1/891 = 0.0011223345
      10'd892: inv_x_count = 16'b0000000001001001; // 1/892 = 0.0011210762
      10'd893: inv_x_count = 16'b0000000001001001; // 1/893 = 0.0011198208
      10'd894: inv_x_count = 16'b0000000001001001; // 1/894 = 0.0011185682
      10'd895: inv_x_count = 16'b0000000001001001; // 1/895 = 0.0011173184
      10'd896: inv_x_count = 16'b0000000001001001; // 1/896 = 0.0011160714
      10'd897: inv_x_count = 16'b0000000001001001; // 1/897 = 0.0011148272
      10'd898: inv_x_count = 16'b0000000001001001; // 1/898 = 0.0011135857
      10'd899: inv_x_count = 16'b0000000001001001; // 1/899 = 0.0011123471
      10'd900: inv_x_count = 16'b0000000001001001; // 1/900 = 0.0011111111
      10'd901: inv_x_count = 16'b0000000001001001; // 1/901 = 0.0011098779
      10'd902: inv_x_count = 16'b0000000001001001; // 1/902 = 0.0011086475
      10'd903: inv_x_count = 16'b0000000001001001; // 1/903 = 0.0011074197
      10'd904: inv_x_count = 16'b0000000001001000; // 1/904 = 0.0011061947
      10'd905: inv_x_count = 16'b0000000001001000; // 1/905 = 0.0011049724
      10'd906: inv_x_count = 16'b0000000001001000; // 1/906 = 0.0011037528
      10'd907: inv_x_count = 16'b0000000001001000; // 1/907 = 0.0011025358
      10'd908: inv_x_count = 16'b0000000001001000; // 1/908 = 0.0011013216
      10'd909: inv_x_count = 16'b0000000001001000; // 1/909 = 0.0011001100
      10'd910: inv_x_count = 16'b0000000001001000; // 1/910 = 0.0010989011
      10'd911: inv_x_count = 16'b0000000001001000; // 1/911 = 0.0010976948
      10'd912: inv_x_count = 16'b0000000001001000; // 1/912 = 0.0010964912
      10'd913: inv_x_count = 16'b0000000001001000; // 1/913 = 0.0010952903
      10'd914: inv_x_count = 16'b0000000001001000; // 1/914 = 0.0010940919
      10'd915: inv_x_count = 16'b0000000001001000; // 1/915 = 0.0010928962
      10'd916: inv_x_count = 16'b0000000001001000; // 1/916 = 0.0010917031
      10'd917: inv_x_count = 16'b0000000001000111; // 1/917 = 0.0010905125
      10'd918: inv_x_count = 16'b0000000001000111; // 1/918 = 0.0010893246
      10'd919: inv_x_count = 16'b0000000001000111; // 1/919 = 0.0010881393
      10'd920: inv_x_count = 16'b0000000001000111; // 1/920 = 0.0010869565
      10'd921: inv_x_count = 16'b0000000001000111; // 1/921 = 0.0010857763
      10'd922: inv_x_count = 16'b0000000001000111; // 1/922 = 0.0010845987
      10'd923: inv_x_count = 16'b0000000001000111; // 1/923 = 0.0010834236
      10'd924: inv_x_count = 16'b0000000001000111; // 1/924 = 0.0010822511
      10'd925: inv_x_count = 16'b0000000001000111; // 1/925 = 0.0010810811
      10'd926: inv_x_count = 16'b0000000001000111; // 1/926 = 0.0010799136
      10'd927: inv_x_count = 16'b0000000001000111; // 1/927 = 0.0010787487
      10'd928: inv_x_count = 16'b0000000001000111; // 1/928 = 0.0010775862
      10'd929: inv_x_count = 16'b0000000001000111; // 1/929 = 0.0010764263
      10'd930: inv_x_count = 16'b0000000001000110; // 1/930 = 0.0010752688
      10'd931: inv_x_count = 16'b0000000001000110; // 1/931 = 0.0010741139
      10'd932: inv_x_count = 16'b0000000001000110; // 1/932 = 0.0010729614
      10'd933: inv_x_count = 16'b0000000001000110; // 1/933 = 0.0010718114
      10'd934: inv_x_count = 16'b0000000001000110; // 1/934 = 0.0010706638
      10'd935: inv_x_count = 16'b0000000001000110; // 1/935 = 0.0010695187
      10'd936: inv_x_count = 16'b0000000001000110; // 1/936 = 0.0010683761
      10'd937: inv_x_count = 16'b0000000001000110; // 1/937 = 0.0010672359
      10'd938: inv_x_count = 16'b0000000001000110; // 1/938 = 0.0010660981
      10'd939: inv_x_count = 16'b0000000001000110; // 1/939 = 0.0010649627
      10'd940: inv_x_count = 16'b0000000001000110; // 1/940 = 0.0010638298
      10'd941: inv_x_count = 16'b0000000001000110; // 1/941 = 0.0010626993
      10'd942: inv_x_count = 16'b0000000001000110; // 1/942 = 0.0010615711
      10'd943: inv_x_count = 16'b0000000001000101; // 1/943 = 0.0010604454
      10'd944: inv_x_count = 16'b0000000001000101; // 1/944 = 0.0010593220
      10'd945: inv_x_count = 16'b0000000001000101; // 1/945 = 0.0010582011
      10'd946: inv_x_count = 16'b0000000001000101; // 1/946 = 0.0010570825
      10'd947: inv_x_count = 16'b0000000001000101; // 1/947 = 0.0010559662
      10'd948: inv_x_count = 16'b0000000001000101; // 1/948 = 0.0010548523
      10'd949: inv_x_count = 16'b0000000001000101; // 1/949 = 0.0010537408
      10'd950: inv_x_count = 16'b0000000001000101; // 1/950 = 0.0010526316
      10'd951: inv_x_count = 16'b0000000001000101; // 1/951 = 0.0010515247
      10'd952: inv_x_count = 16'b0000000001000101; // 1/952 = 0.0010504202
      10'd953: inv_x_count = 16'b0000000001000101; // 1/953 = 0.0010493179
      10'd954: inv_x_count = 16'b0000000001000101; // 1/954 = 0.0010482180
      10'd955: inv_x_count = 16'b0000000001000101; // 1/955 = 0.0010471204
      10'd956: inv_x_count = 16'b0000000001000101; // 1/956 = 0.0010460251
      10'd957: inv_x_count = 16'b0000000001000100; // 1/957 = 0.0010449321
      10'd958: inv_x_count = 16'b0000000001000100; // 1/958 = 0.0010438413
      10'd959: inv_x_count = 16'b0000000001000100; // 1/959 = 0.0010427529
      10'd960: inv_x_count = 16'b0000000001000100; // 1/960 = 0.0010416667
      10'd961: inv_x_count = 16'b0000000001000100; // 1/961 = 0.0010405827
      10'd962: inv_x_count = 16'b0000000001000100; // 1/962 = 0.0010395010
      10'd963: inv_x_count = 16'b0000000001000100; // 1/963 = 0.0010384216
      10'd964: inv_x_count = 16'b0000000001000100; // 1/964 = 0.0010373444
      10'd965: inv_x_count = 16'b0000000001000100; // 1/965 = 0.0010362694
      10'd966: inv_x_count = 16'b0000000001000100; // 1/966 = 0.0010351967
      10'd967: inv_x_count = 16'b0000000001000100; // 1/967 = 0.0010341262
      10'd968: inv_x_count = 16'b0000000001000100; // 1/968 = 0.0010330579
      10'd969: inv_x_count = 16'b0000000001000100; // 1/969 = 0.0010319917
      10'd970: inv_x_count = 16'b0000000001000100; // 1/970 = 0.0010309278
      10'd971: inv_x_count = 16'b0000000001000011; // 1/971 = 0.0010298661
      10'd972: inv_x_count = 16'b0000000001000011; // 1/972 = 0.0010288066
      10'd973: inv_x_count = 16'b0000000001000011; // 1/973 = 0.0010277492
      10'd974: inv_x_count = 16'b0000000001000011; // 1/974 = 0.0010266940
      10'd975: inv_x_count = 16'b0000000001000011; // 1/975 = 0.0010256410
      10'd976: inv_x_count = 16'b0000000001000011; // 1/976 = 0.0010245902
      10'd977: inv_x_count = 16'b0000000001000011; // 1/977 = 0.0010235415
      10'd978: inv_x_count = 16'b0000000001000011; // 1/978 = 0.0010224949
      10'd979: inv_x_count = 16'b0000000001000011; // 1/979 = 0.0010214505
      10'd980: inv_x_count = 16'b0000000001000011; // 1/980 = 0.0010204082
      10'd981: inv_x_count = 16'b0000000001000011; // 1/981 = 0.0010193680
      10'd982: inv_x_count = 16'b0000000001000011; // 1/982 = 0.0010183299
      10'd983: inv_x_count = 16'b0000000001000011; // 1/983 = 0.0010172940
      10'd984: inv_x_count = 16'b0000000001000011; // 1/984 = 0.0010162602
      10'd985: inv_x_count = 16'b0000000001000011; // 1/985 = 0.0010152284
      10'd986: inv_x_count = 16'b0000000001000010; // 1/986 = 0.0010141988
      10'd987: inv_x_count = 16'b0000000001000010; // 1/987 = 0.0010131712
      10'd988: inv_x_count = 16'b0000000001000010; // 1/988 = 0.0010121457
      10'd989: inv_x_count = 16'b0000000001000010; // 1/989 = 0.0010111223
      10'd990: inv_x_count = 16'b0000000001000010; // 1/990 = 0.0010101010
      10'd991: inv_x_count = 16'b0000000001000010; // 1/991 = 0.0010090817
      10'd992: inv_x_count = 16'b0000000001000010; // 1/992 = 0.0010080645
      10'd993: inv_x_count = 16'b0000000001000010; // 1/993 = 0.0010070493
      10'd994: inv_x_count = 16'b0000000001000010; // 1/994 = 0.0010060362
      10'd995: inv_x_count = 16'b0000000001000010; // 1/995 = 0.0010050251
      10'd996: inv_x_count = 16'b0000000001000010; // 1/996 = 0.0010040161
      10'd997: inv_x_count = 16'b0000000001000010; // 1/997 = 0.0010030090
      10'd998: inv_x_count = 16'b0000000001000010; // 1/998 = 0.0010020040
      10'd999: inv_x_count = 16'b0000000001000010; // 1/999 = 0.0010010010
      10'd1000: inv_x_count = 16'b0000000001000010; // 1/1000 = 0.0010000000
      10'd1001: inv_x_count = 16'b0000000001000001; // 1/1001 = 0.0009990010
      10'd1002: inv_x_count = 16'b0000000001000001; // 1/1002 = 0.0009980040
      10'd1003: inv_x_count = 16'b0000000001000001; // 1/1003 = 0.0009970090
      10'd1004: inv_x_count = 16'b0000000001000001; // 1/1004 = 0.0009960159
      10'd1005: inv_x_count = 16'b0000000001000001; // 1/1005 = 0.0009950249
      10'd1006: inv_x_count = 16'b0000000001000001; // 1/1006 = 0.0009940358
      10'd1007: inv_x_count = 16'b0000000001000001; // 1/1007 = 0.0009930487
      10'd1008: inv_x_count = 16'b0000000001000001; // 1/1008 = 0.0009920635
      10'd1009: inv_x_count = 16'b0000000001000001; // 1/1009 = 0.0009910803
      10'd1010: inv_x_count = 16'b0000000001000001; // 1/1010 = 0.0009900990
      10'd1011: inv_x_count = 16'b0000000001000001; // 1/1011 = 0.0009891197
      10'd1012: inv_x_count = 16'b0000000001000001; // 1/1012 = 0.0009881423
      10'd1013: inv_x_count = 16'b0000000001000001; // 1/1013 = 0.0009871668
      10'd1014: inv_x_count = 16'b0000000001000001; // 1/1014 = 0.0009861933
      10'd1015: inv_x_count = 16'b0000000001000001; // 1/1015 = 0.0009852217
      10'd1016: inv_x_count = 16'b0000000001000001; // 1/1016 = 0.0009842520
      10'd1017: inv_x_count = 16'b0000000001000000; // 1/1017 = 0.0009832842
      10'd1018: inv_x_count = 16'b0000000001000000; // 1/1018 = 0.0009823183
      10'd1019: inv_x_count = 16'b0000000001000000; // 1/1019 = 0.0009813543
      10'd1020: inv_x_count = 16'b0000000001000000; // 1/1020 = 0.0009803922
      10'd1021: inv_x_count = 16'b0000000001000000; // 1/1021 = 0.0009794319
      10'd1022: inv_x_count = 16'b0000000001000000; // 1/1022 = 0.0009784736
      10'd1023: inv_x_count = 16'b0000000001000000; // 1/1023 = 0.0009775171
      10'd1024: inv_x_count = 16'b0000000001000000; // 1/1024 = 0.0009765625
      default: inv_x_count = '0; // Default case
    endcase
  end

  always_comb begin
    case (x_count-1)
      10'd2: inv_x_count_prev = 16'b1000000000000000; // 1/2 = 0.5000000000
      10'd3: inv_x_count_prev = 16'b0101010101010101; // 1/3 = 0.3333333333
      10'd4: inv_x_count_prev = 16'b0100000000000000; // 1/4 = 0.2500000000
      10'd5: inv_x_count_prev = 16'b0011001100110011; // 1/5 = 0.2000000000
      10'd6: inv_x_count_prev = 16'b0010101010101011; // 1/6 = 0.1666666667
      10'd7: inv_x_count_prev = 16'b0010010010010010; // 1/7 = 0.1428571429
      10'd8: inv_x_count_prev = 16'b0010000000000000; // 1/8 = 0.1250000000
      10'd9: inv_x_count_prev = 16'b0001110001110010; // 1/9 = 0.1111111111
      10'd10: inv_x_count_prev = 16'b0001100110011010; // 1/10 = 0.1000000000
      10'd11: inv_x_count_prev = 16'b0001011101000110; // 1/11 = 0.0909090909
      10'd12: inv_x_count_prev = 16'b0001010101010101; // 1/12 = 0.0833333333
      10'd13: inv_x_count_prev = 16'b0001001110110001; // 1/13 = 0.0769230769
      10'd14: inv_x_count_prev = 16'b0001001001001001; // 1/14 = 0.0714285714
      10'd15: inv_x_count_prev = 16'b0001000100010001; // 1/15 = 0.0666666667
      10'd16: inv_x_count_prev = 16'b0001000000000000; // 1/16 = 0.0625000000
      10'd17: inv_x_count_prev = 16'b0000111100001111; // 1/17 = 0.0588235294
      10'd18: inv_x_count_prev = 16'b0000111000111001; // 1/18 = 0.0555555556
      10'd19: inv_x_count_prev = 16'b0000110101111001; // 1/19 = 0.0526315789
      10'd20: inv_x_count_prev = 16'b0000110011001101; // 1/20 = 0.0500000000
      10'd21: inv_x_count_prev = 16'b0000110000110001; // 1/21 = 0.0476190476
      10'd22: inv_x_count_prev = 16'b0000101110100011; // 1/22 = 0.0454545455
      10'd23: inv_x_count_prev = 16'b0000101100100001; // 1/23 = 0.0434782609
      10'd24: inv_x_count_prev = 16'b0000101010101011; // 1/24 = 0.0416666667
      10'd25: inv_x_count_prev = 16'b0000101000111101; // 1/25 = 0.0400000000
      10'd26: inv_x_count_prev = 16'b0000100111011001; // 1/26 = 0.0384615385
      10'd27: inv_x_count_prev = 16'b0000100101111011; // 1/27 = 0.0370370370
      10'd28: inv_x_count_prev = 16'b0000100100100101; // 1/28 = 0.0357142857
      10'd29: inv_x_count_prev = 16'b0000100011010100; // 1/29 = 0.0344827586
      10'd30: inv_x_count_prev = 16'b0000100010001001; // 1/30 = 0.0333333333
      10'd31: inv_x_count_prev = 16'b0000100001000010; // 1/31 = 0.0322580645
      10'd32: inv_x_count_prev = 16'b0000100000000000; // 1/32 = 0.0312500000
      10'd33: inv_x_count_prev = 16'b0000011111000010; // 1/33 = 0.0303030303
      10'd34: inv_x_count_prev = 16'b0000011110001000; // 1/34 = 0.0294117647
      10'd35: inv_x_count_prev = 16'b0000011101010000; // 1/35 = 0.0285714286
      10'd36: inv_x_count_prev = 16'b0000011100011100; // 1/36 = 0.0277777778
      10'd37: inv_x_count_prev = 16'b0000011011101011; // 1/37 = 0.0270270270
      10'd38: inv_x_count_prev = 16'b0000011010111101; // 1/38 = 0.0263157895
      10'd39: inv_x_count_prev = 16'b0000011010010000; // 1/39 = 0.0256410256
      10'd40: inv_x_count_prev = 16'b0000011001100110; // 1/40 = 0.0250000000
      10'd41: inv_x_count_prev = 16'b0000011000111110; // 1/41 = 0.0243902439
      10'd42: inv_x_count_prev = 16'b0000011000011000; // 1/42 = 0.0238095238
      10'd43: inv_x_count_prev = 16'b0000010111110100; // 1/43 = 0.0232558140
      10'd44: inv_x_count_prev = 16'b0000010111010001; // 1/44 = 0.0227272727
      10'd45: inv_x_count_prev = 16'b0000010110110000; // 1/45 = 0.0222222222
      10'd46: inv_x_count_prev = 16'b0000010110010001; // 1/46 = 0.0217391304
      10'd47: inv_x_count_prev = 16'b0000010101110010; // 1/47 = 0.0212765957
      10'd48: inv_x_count_prev = 16'b0000010101010101; // 1/48 = 0.0208333333
      10'd49: inv_x_count_prev = 16'b0000010100111001; // 1/49 = 0.0204081633
      10'd50: inv_x_count_prev = 16'b0000010100011111; // 1/50 = 0.0200000000
      10'd51: inv_x_count_prev = 16'b0000010100000101; // 1/51 = 0.0196078431
      10'd52: inv_x_count_prev = 16'b0000010011101100; // 1/52 = 0.0192307692
      10'd53: inv_x_count_prev = 16'b0000010011010101; // 1/53 = 0.0188679245
      10'd54: inv_x_count_prev = 16'b0000010010111110; // 1/54 = 0.0185185185
      10'd55: inv_x_count_prev = 16'b0000010010101000; // 1/55 = 0.0181818182
      10'd56: inv_x_count_prev = 16'b0000010010010010; // 1/56 = 0.0178571429
      10'd57: inv_x_count_prev = 16'b0000010001111110; // 1/57 = 0.0175438596
      10'd58: inv_x_count_prev = 16'b0000010001101010; // 1/58 = 0.0172413793
      10'd59: inv_x_count_prev = 16'b0000010001010111; // 1/59 = 0.0169491525
      10'd60: inv_x_count_prev = 16'b0000010001000100; // 1/60 = 0.0166666667
      10'd61: inv_x_count_prev = 16'b0000010000110010; // 1/61 = 0.0163934426
      10'd62: inv_x_count_prev = 16'b0000010000100001; // 1/62 = 0.0161290323
      10'd63: inv_x_count_prev = 16'b0000010000010000; // 1/63 = 0.0158730159
      10'd64: inv_x_count_prev = 16'b0000010000000000; // 1/64 = 0.0156250000
      10'd65: inv_x_count_prev = 16'b0000001111110000; // 1/65 = 0.0153846154
      10'd66: inv_x_count_prev = 16'b0000001111100001; // 1/66 = 0.0151515152
      10'd67: inv_x_count_prev = 16'b0000001111010010; // 1/67 = 0.0149253731
      10'd68: inv_x_count_prev = 16'b0000001111000100; // 1/68 = 0.0147058824
      10'd69: inv_x_count_prev = 16'b0000001110110110; // 1/69 = 0.0144927536
      10'd70: inv_x_count_prev = 16'b0000001110101000; // 1/70 = 0.0142857143
      10'd71: inv_x_count_prev = 16'b0000001110011011; // 1/71 = 0.0140845070
      10'd72: inv_x_count_prev = 16'b0000001110001110; // 1/72 = 0.0138888889
      10'd73: inv_x_count_prev = 16'b0000001110000010; // 1/73 = 0.0136986301
      10'd74: inv_x_count_prev = 16'b0000001101110110; // 1/74 = 0.0135135135
      10'd75: inv_x_count_prev = 16'b0000001101101010; // 1/75 = 0.0133333333
      10'd76: inv_x_count_prev = 16'b0000001101011110; // 1/76 = 0.0131578947
      10'd77: inv_x_count_prev = 16'b0000001101010011; // 1/77 = 0.0129870130
      10'd78: inv_x_count_prev = 16'b0000001101001000; // 1/78 = 0.0128205128
      10'd79: inv_x_count_prev = 16'b0000001100111110; // 1/79 = 0.0126582278
      10'd80: inv_x_count_prev = 16'b0000001100110011; // 1/80 = 0.0125000000
      10'd81: inv_x_count_prev = 16'b0000001100101001; // 1/81 = 0.0123456790
      10'd82: inv_x_count_prev = 16'b0000001100011111; // 1/82 = 0.0121951220
      10'd83: inv_x_count_prev = 16'b0000001100010110; // 1/83 = 0.0120481928
      10'd84: inv_x_count_prev = 16'b0000001100001100; // 1/84 = 0.0119047619
      10'd85: inv_x_count_prev = 16'b0000001100000011; // 1/85 = 0.0117647059
      10'd86: inv_x_count_prev = 16'b0000001011111010; // 1/86 = 0.0116279070
      10'd87: inv_x_count_prev = 16'b0000001011110001; // 1/87 = 0.0114942529
      10'd88: inv_x_count_prev = 16'b0000001011101001; // 1/88 = 0.0113636364
      10'd89: inv_x_count_prev = 16'b0000001011100000; // 1/89 = 0.0112359551
      10'd90: inv_x_count_prev = 16'b0000001011011000; // 1/90 = 0.0111111111
      10'd91: inv_x_count_prev = 16'b0000001011010000; // 1/91 = 0.0109890110
      10'd92: inv_x_count_prev = 16'b0000001011001000; // 1/92 = 0.0108695652
      10'd93: inv_x_count_prev = 16'b0000001011000001; // 1/93 = 0.0107526882
      10'd94: inv_x_count_prev = 16'b0000001010111001; // 1/94 = 0.0106382979
      10'd95: inv_x_count_prev = 16'b0000001010110010; // 1/95 = 0.0105263158
      10'd96: inv_x_count_prev = 16'b0000001010101011; // 1/96 = 0.0104166667
      10'd97: inv_x_count_prev = 16'b0000001010100100; // 1/97 = 0.0103092784
      10'd98: inv_x_count_prev = 16'b0000001010011101; // 1/98 = 0.0102040816
      10'd99: inv_x_count_prev = 16'b0000001010010110; // 1/99 = 0.0101010101
      10'd100: inv_x_count_prev = 16'b0000001010001111; // 1/100 = 0.0100000000
      10'd101: inv_x_count_prev = 16'b0000001010001001; // 1/101 = 0.0099009901
      10'd102: inv_x_count_prev = 16'b0000001010000011; // 1/102 = 0.0098039216
      10'd103: inv_x_count_prev = 16'b0000001001111100; // 1/103 = 0.0097087379
      10'd104: inv_x_count_prev = 16'b0000001001110110; // 1/104 = 0.0096153846
      10'd105: inv_x_count_prev = 16'b0000001001110000; // 1/105 = 0.0095238095
      10'd106: inv_x_count_prev = 16'b0000001001101010; // 1/106 = 0.0094339623
      10'd107: inv_x_count_prev = 16'b0000001001100100; // 1/107 = 0.0093457944
      10'd108: inv_x_count_prev = 16'b0000001001011111; // 1/108 = 0.0092592593
      10'd109: inv_x_count_prev = 16'b0000001001011001; // 1/109 = 0.0091743119
      10'd110: inv_x_count_prev = 16'b0000001001010100; // 1/110 = 0.0090909091
      10'd111: inv_x_count_prev = 16'b0000001001001110; // 1/111 = 0.0090090090
      10'd112: inv_x_count_prev = 16'b0000001001001001; // 1/112 = 0.0089285714
      10'd113: inv_x_count_prev = 16'b0000001001000100; // 1/113 = 0.0088495575
      10'd114: inv_x_count_prev = 16'b0000001000111111; // 1/114 = 0.0087719298
      10'd115: inv_x_count_prev = 16'b0000001000111010; // 1/115 = 0.0086956522
      10'd116: inv_x_count_prev = 16'b0000001000110101; // 1/116 = 0.0086206897
      10'd117: inv_x_count_prev = 16'b0000001000110000; // 1/117 = 0.0085470085
      10'd118: inv_x_count_prev = 16'b0000001000101011; // 1/118 = 0.0084745763
      10'd119: inv_x_count_prev = 16'b0000001000100111; // 1/119 = 0.0084033613
      10'd120: inv_x_count_prev = 16'b0000001000100010; // 1/120 = 0.0083333333
      10'd121: inv_x_count_prev = 16'b0000001000011110; // 1/121 = 0.0082644628
      10'd122: inv_x_count_prev = 16'b0000001000011001; // 1/122 = 0.0081967213
      10'd123: inv_x_count_prev = 16'b0000001000010101; // 1/123 = 0.0081300813
      10'd124: inv_x_count_prev = 16'b0000001000010001; // 1/124 = 0.0080645161
      10'd125: inv_x_count_prev = 16'b0000001000001100; // 1/125 = 0.0080000000
      10'd126: inv_x_count_prev = 16'b0000001000001000; // 1/126 = 0.0079365079
      10'd127: inv_x_count_prev = 16'b0000001000000100; // 1/127 = 0.0078740157
      10'd128: inv_x_count_prev = 16'b0000001000000000; // 1/128 = 0.0078125000
      10'd129: inv_x_count_prev = 16'b0000000111111100; // 1/129 = 0.0077519380
      10'd130: inv_x_count_prev = 16'b0000000111111000; // 1/130 = 0.0076923077
      10'd131: inv_x_count_prev = 16'b0000000111110100; // 1/131 = 0.0076335878
      10'd132: inv_x_count_prev = 16'b0000000111110000; // 1/132 = 0.0075757576
      10'd133: inv_x_count_prev = 16'b0000000111101101; // 1/133 = 0.0075187970
      10'd134: inv_x_count_prev = 16'b0000000111101001; // 1/134 = 0.0074626866
      10'd135: inv_x_count_prev = 16'b0000000111100101; // 1/135 = 0.0074074074
      10'd136: inv_x_count_prev = 16'b0000000111100010; // 1/136 = 0.0073529412
      10'd137: inv_x_count_prev = 16'b0000000111011110; // 1/137 = 0.0072992701
      10'd138: inv_x_count_prev = 16'b0000000111011011; // 1/138 = 0.0072463768
      10'd139: inv_x_count_prev = 16'b0000000111010111; // 1/139 = 0.0071942446
      10'd140: inv_x_count_prev = 16'b0000000111010100; // 1/140 = 0.0071428571
      10'd141: inv_x_count_prev = 16'b0000000111010001; // 1/141 = 0.0070921986
      10'd142: inv_x_count_prev = 16'b0000000111001110; // 1/142 = 0.0070422535
      10'd143: inv_x_count_prev = 16'b0000000111001010; // 1/143 = 0.0069930070
      10'd144: inv_x_count_prev = 16'b0000000111000111; // 1/144 = 0.0069444444
      10'd145: inv_x_count_prev = 16'b0000000111000100; // 1/145 = 0.0068965517
      10'd146: inv_x_count_prev = 16'b0000000111000001; // 1/146 = 0.0068493151
      10'd147: inv_x_count_prev = 16'b0000000110111110; // 1/147 = 0.0068027211
      10'd148: inv_x_count_prev = 16'b0000000110111011; // 1/148 = 0.0067567568
      10'd149: inv_x_count_prev = 16'b0000000110111000; // 1/149 = 0.0067114094
      10'd150: inv_x_count_prev = 16'b0000000110110101; // 1/150 = 0.0066666667
      10'd151: inv_x_count_prev = 16'b0000000110110010; // 1/151 = 0.0066225166
      10'd152: inv_x_count_prev = 16'b0000000110101111; // 1/152 = 0.0065789474
      10'd153: inv_x_count_prev = 16'b0000000110101100; // 1/153 = 0.0065359477
      10'd154: inv_x_count_prev = 16'b0000000110101010; // 1/154 = 0.0064935065
      10'd155: inv_x_count_prev = 16'b0000000110100111; // 1/155 = 0.0064516129
      10'd156: inv_x_count_prev = 16'b0000000110100100; // 1/156 = 0.0064102564
      10'd157: inv_x_count_prev = 16'b0000000110100001; // 1/157 = 0.0063694268
      10'd158: inv_x_count_prev = 16'b0000000110011111; // 1/158 = 0.0063291139
      10'd159: inv_x_count_prev = 16'b0000000110011100; // 1/159 = 0.0062893082
      10'd160: inv_x_count_prev = 16'b0000000110011010; // 1/160 = 0.0062500000
      10'd161: inv_x_count_prev = 16'b0000000110010111; // 1/161 = 0.0062111801
      10'd162: inv_x_count_prev = 16'b0000000110010101; // 1/162 = 0.0061728395
      10'd163: inv_x_count_prev = 16'b0000000110010010; // 1/163 = 0.0061349693
      10'd164: inv_x_count_prev = 16'b0000000110010000; // 1/164 = 0.0060975610
      10'd165: inv_x_count_prev = 16'b0000000110001101; // 1/165 = 0.0060606061
      10'd166: inv_x_count_prev = 16'b0000000110001011; // 1/166 = 0.0060240964
      10'd167: inv_x_count_prev = 16'b0000000110001000; // 1/167 = 0.0059880240
      10'd168: inv_x_count_prev = 16'b0000000110000110; // 1/168 = 0.0059523810
      10'd169: inv_x_count_prev = 16'b0000000110000100; // 1/169 = 0.0059171598
      10'd170: inv_x_count_prev = 16'b0000000110000010; // 1/170 = 0.0058823529
      10'd171: inv_x_count_prev = 16'b0000000101111111; // 1/171 = 0.0058479532
      10'd172: inv_x_count_prev = 16'b0000000101111101; // 1/172 = 0.0058139535
      10'd173: inv_x_count_prev = 16'b0000000101111011; // 1/173 = 0.0057803468
      10'd174: inv_x_count_prev = 16'b0000000101111001; // 1/174 = 0.0057471264
      10'd175: inv_x_count_prev = 16'b0000000101110110; // 1/175 = 0.0057142857
      10'd176: inv_x_count_prev = 16'b0000000101110100; // 1/176 = 0.0056818182
      10'd177: inv_x_count_prev = 16'b0000000101110010; // 1/177 = 0.0056497175
      10'd178: inv_x_count_prev = 16'b0000000101110000; // 1/178 = 0.0056179775
      10'd179: inv_x_count_prev = 16'b0000000101101110; // 1/179 = 0.0055865922
      10'd180: inv_x_count_prev = 16'b0000000101101100; // 1/180 = 0.0055555556
      10'd181: inv_x_count_prev = 16'b0000000101101010; // 1/181 = 0.0055248619
      10'd182: inv_x_count_prev = 16'b0000000101101000; // 1/182 = 0.0054945055
      10'd183: inv_x_count_prev = 16'b0000000101100110; // 1/183 = 0.0054644809
      10'd184: inv_x_count_prev = 16'b0000000101100100; // 1/184 = 0.0054347826
      10'd185: inv_x_count_prev = 16'b0000000101100010; // 1/185 = 0.0054054054
      10'd186: inv_x_count_prev = 16'b0000000101100000; // 1/186 = 0.0053763441
      10'd187: inv_x_count_prev = 16'b0000000101011110; // 1/187 = 0.0053475936
      10'd188: inv_x_count_prev = 16'b0000000101011101; // 1/188 = 0.0053191489
      10'd189: inv_x_count_prev = 16'b0000000101011011; // 1/189 = 0.0052910053
      10'd190: inv_x_count_prev = 16'b0000000101011001; // 1/190 = 0.0052631579
      10'd191: inv_x_count_prev = 16'b0000000101010111; // 1/191 = 0.0052356021
      10'd192: inv_x_count_prev = 16'b0000000101010101; // 1/192 = 0.0052083333
      10'd193: inv_x_count_prev = 16'b0000000101010100; // 1/193 = 0.0051813472
      10'd194: inv_x_count_prev = 16'b0000000101010010; // 1/194 = 0.0051546392
      10'd195: inv_x_count_prev = 16'b0000000101010000; // 1/195 = 0.0051282051
      10'd196: inv_x_count_prev = 16'b0000000101001110; // 1/196 = 0.0051020408
      10'd197: inv_x_count_prev = 16'b0000000101001101; // 1/197 = 0.0050761421
      10'd198: inv_x_count_prev = 16'b0000000101001011; // 1/198 = 0.0050505051
      10'd199: inv_x_count_prev = 16'b0000000101001001; // 1/199 = 0.0050251256
      10'd200: inv_x_count_prev = 16'b0000000101001000; // 1/200 = 0.0050000000
      10'd201: inv_x_count_prev = 16'b0000000101000110; // 1/201 = 0.0049751244
      10'd202: inv_x_count_prev = 16'b0000000101000100; // 1/202 = 0.0049504950
      10'd203: inv_x_count_prev = 16'b0000000101000011; // 1/203 = 0.0049261084
      10'd204: inv_x_count_prev = 16'b0000000101000001; // 1/204 = 0.0049019608
      10'd205: inv_x_count_prev = 16'b0000000101000000; // 1/205 = 0.0048780488
      10'd206: inv_x_count_prev = 16'b0000000100111110; // 1/206 = 0.0048543689
      10'd207: inv_x_count_prev = 16'b0000000100111101; // 1/207 = 0.0048309179
      10'd208: inv_x_count_prev = 16'b0000000100111011; // 1/208 = 0.0048076923
      10'd209: inv_x_count_prev = 16'b0000000100111010; // 1/209 = 0.0047846890
      10'd210: inv_x_count_prev = 16'b0000000100111000; // 1/210 = 0.0047619048
      10'd211: inv_x_count_prev = 16'b0000000100110111; // 1/211 = 0.0047393365
      10'd212: inv_x_count_prev = 16'b0000000100110101; // 1/212 = 0.0047169811
      10'd213: inv_x_count_prev = 16'b0000000100110100; // 1/213 = 0.0046948357
      10'd214: inv_x_count_prev = 16'b0000000100110010; // 1/214 = 0.0046728972
      10'd215: inv_x_count_prev = 16'b0000000100110001; // 1/215 = 0.0046511628
      10'd216: inv_x_count_prev = 16'b0000000100101111; // 1/216 = 0.0046296296
      10'd217: inv_x_count_prev = 16'b0000000100101110; // 1/217 = 0.0046082949
      10'd218: inv_x_count_prev = 16'b0000000100101101; // 1/218 = 0.0045871560
      10'd219: inv_x_count_prev = 16'b0000000100101011; // 1/219 = 0.0045662100
      10'd220: inv_x_count_prev = 16'b0000000100101010; // 1/220 = 0.0045454545
      10'd221: inv_x_count_prev = 16'b0000000100101001; // 1/221 = 0.0045248869
      10'd222: inv_x_count_prev = 16'b0000000100100111; // 1/222 = 0.0045045045
      10'd223: inv_x_count_prev = 16'b0000000100100110; // 1/223 = 0.0044843049
      10'd224: inv_x_count_prev = 16'b0000000100100101; // 1/224 = 0.0044642857
      10'd225: inv_x_count_prev = 16'b0000000100100011; // 1/225 = 0.0044444444
      10'd226: inv_x_count_prev = 16'b0000000100100010; // 1/226 = 0.0044247788
      10'd227: inv_x_count_prev = 16'b0000000100100001; // 1/227 = 0.0044052863
      10'd228: inv_x_count_prev = 16'b0000000100011111; // 1/228 = 0.0043859649
      10'd229: inv_x_count_prev = 16'b0000000100011110; // 1/229 = 0.0043668122
      10'd230: inv_x_count_prev = 16'b0000000100011101; // 1/230 = 0.0043478261
      10'd231: inv_x_count_prev = 16'b0000000100011100; // 1/231 = 0.0043290043
      10'd232: inv_x_count_prev = 16'b0000000100011010; // 1/232 = 0.0043103448
      10'd233: inv_x_count_prev = 16'b0000000100011001; // 1/233 = 0.0042918455
      10'd234: inv_x_count_prev = 16'b0000000100011000; // 1/234 = 0.0042735043
      10'd235: inv_x_count_prev = 16'b0000000100010111; // 1/235 = 0.0042553191
      10'd236: inv_x_count_prev = 16'b0000000100010110; // 1/236 = 0.0042372881
      10'd237: inv_x_count_prev = 16'b0000000100010101; // 1/237 = 0.0042194093
      10'd238: inv_x_count_prev = 16'b0000000100010011; // 1/238 = 0.0042016807
      10'd239: inv_x_count_prev = 16'b0000000100010010; // 1/239 = 0.0041841004
      10'd240: inv_x_count_prev = 16'b0000000100010001; // 1/240 = 0.0041666667
      10'd241: inv_x_count_prev = 16'b0000000100010000; // 1/241 = 0.0041493776
      10'd242: inv_x_count_prev = 16'b0000000100001111; // 1/242 = 0.0041322314
      10'd243: inv_x_count_prev = 16'b0000000100001110; // 1/243 = 0.0041152263
      10'd244: inv_x_count_prev = 16'b0000000100001101; // 1/244 = 0.0040983607
      10'd245: inv_x_count_prev = 16'b0000000100001011; // 1/245 = 0.0040816327
      10'd246: inv_x_count_prev = 16'b0000000100001010; // 1/246 = 0.0040650407
      10'd247: inv_x_count_prev = 16'b0000000100001001; // 1/247 = 0.0040485830
      10'd248: inv_x_count_prev = 16'b0000000100001000; // 1/248 = 0.0040322581
      10'd249: inv_x_count_prev = 16'b0000000100000111; // 1/249 = 0.0040160643
      10'd250: inv_x_count_prev = 16'b0000000100000110; // 1/250 = 0.0040000000
      10'd251: inv_x_count_prev = 16'b0000000100000101; // 1/251 = 0.0039840637
      10'd252: inv_x_count_prev = 16'b0000000100000100; // 1/252 = 0.0039682540
      10'd253: inv_x_count_prev = 16'b0000000100000011; // 1/253 = 0.0039525692
      10'd254: inv_x_count_prev = 16'b0000000100000010; // 1/254 = 0.0039370079
      10'd255: inv_x_count_prev = 16'b0000000100000001; // 1/255 = 0.0039215686
      10'd256: inv_x_count_prev = 16'b0000000100000000; // 1/256 = 0.0039062500
      10'd257: inv_x_count_prev = 16'b0000000011111111; // 1/257 = 0.0038910506
      10'd258: inv_x_count_prev = 16'b0000000011111110; // 1/258 = 0.0038759690
      10'd259: inv_x_count_prev = 16'b0000000011111101; // 1/259 = 0.0038610039
      10'd260: inv_x_count_prev = 16'b0000000011111100; // 1/260 = 0.0038461538
      10'd261: inv_x_count_prev = 16'b0000000011111011; // 1/261 = 0.0038314176
      10'd262: inv_x_count_prev = 16'b0000000011111010; // 1/262 = 0.0038167939
      10'd263: inv_x_count_prev = 16'b0000000011111001; // 1/263 = 0.0038022814
      10'd264: inv_x_count_prev = 16'b0000000011111000; // 1/264 = 0.0037878788
      10'd265: inv_x_count_prev = 16'b0000000011110111; // 1/265 = 0.0037735849
      10'd266: inv_x_count_prev = 16'b0000000011110110; // 1/266 = 0.0037593985
      10'd267: inv_x_count_prev = 16'b0000000011110101; // 1/267 = 0.0037453184
      10'd268: inv_x_count_prev = 16'b0000000011110101; // 1/268 = 0.0037313433
      10'd269: inv_x_count_prev = 16'b0000000011110100; // 1/269 = 0.0037174721
      10'd270: inv_x_count_prev = 16'b0000000011110011; // 1/270 = 0.0037037037
      10'd271: inv_x_count_prev = 16'b0000000011110010; // 1/271 = 0.0036900369
      10'd272: inv_x_count_prev = 16'b0000000011110001; // 1/272 = 0.0036764706
      10'd273: inv_x_count_prev = 16'b0000000011110000; // 1/273 = 0.0036630037
      10'd274: inv_x_count_prev = 16'b0000000011101111; // 1/274 = 0.0036496350
      10'd275: inv_x_count_prev = 16'b0000000011101110; // 1/275 = 0.0036363636
      10'd276: inv_x_count_prev = 16'b0000000011101101; // 1/276 = 0.0036231884
      10'd277: inv_x_count_prev = 16'b0000000011101101; // 1/277 = 0.0036101083
      10'd278: inv_x_count_prev = 16'b0000000011101100; // 1/278 = 0.0035971223
      10'd279: inv_x_count_prev = 16'b0000000011101011; // 1/279 = 0.0035842294
      10'd280: inv_x_count_prev = 16'b0000000011101010; // 1/280 = 0.0035714286
      10'd281: inv_x_count_prev = 16'b0000000011101001; // 1/281 = 0.0035587189
      10'd282: inv_x_count_prev = 16'b0000000011101000; // 1/282 = 0.0035460993
      10'd283: inv_x_count_prev = 16'b0000000011101000; // 1/283 = 0.0035335689
      10'd284: inv_x_count_prev = 16'b0000000011100111; // 1/284 = 0.0035211268
      10'd285: inv_x_count_prev = 16'b0000000011100110; // 1/285 = 0.0035087719
      10'd286: inv_x_count_prev = 16'b0000000011100101; // 1/286 = 0.0034965035
      10'd287: inv_x_count_prev = 16'b0000000011100100; // 1/287 = 0.0034843206
      10'd288: inv_x_count_prev = 16'b0000000011100100; // 1/288 = 0.0034722222
      10'd289: inv_x_count_prev = 16'b0000000011100011; // 1/289 = 0.0034602076
      10'd290: inv_x_count_prev = 16'b0000000011100010; // 1/290 = 0.0034482759
      10'd291: inv_x_count_prev = 16'b0000000011100001; // 1/291 = 0.0034364261
      10'd292: inv_x_count_prev = 16'b0000000011100000; // 1/292 = 0.0034246575
      10'd293: inv_x_count_prev = 16'b0000000011100000; // 1/293 = 0.0034129693
      10'd294: inv_x_count_prev = 16'b0000000011011111; // 1/294 = 0.0034013605
      10'd295: inv_x_count_prev = 16'b0000000011011110; // 1/295 = 0.0033898305
      10'd296: inv_x_count_prev = 16'b0000000011011101; // 1/296 = 0.0033783784
      10'd297: inv_x_count_prev = 16'b0000000011011101; // 1/297 = 0.0033670034
      10'd298: inv_x_count_prev = 16'b0000000011011100; // 1/298 = 0.0033557047
      10'd299: inv_x_count_prev = 16'b0000000011011011; // 1/299 = 0.0033444816
      10'd300: inv_x_count_prev = 16'b0000000011011010; // 1/300 = 0.0033333333
      10'd301: inv_x_count_prev = 16'b0000000011011010; // 1/301 = 0.0033222591
      10'd302: inv_x_count_prev = 16'b0000000011011001; // 1/302 = 0.0033112583
      10'd303: inv_x_count_prev = 16'b0000000011011000; // 1/303 = 0.0033003300
      10'd304: inv_x_count_prev = 16'b0000000011011000; // 1/304 = 0.0032894737
      10'd305: inv_x_count_prev = 16'b0000000011010111; // 1/305 = 0.0032786885
      10'd306: inv_x_count_prev = 16'b0000000011010110; // 1/306 = 0.0032679739
      10'd307: inv_x_count_prev = 16'b0000000011010101; // 1/307 = 0.0032573290
      10'd308: inv_x_count_prev = 16'b0000000011010101; // 1/308 = 0.0032467532
      10'd309: inv_x_count_prev = 16'b0000000011010100; // 1/309 = 0.0032362460
      10'd310: inv_x_count_prev = 16'b0000000011010011; // 1/310 = 0.0032258065
      10'd311: inv_x_count_prev = 16'b0000000011010011; // 1/311 = 0.0032154341
      10'd312: inv_x_count_prev = 16'b0000000011010010; // 1/312 = 0.0032051282
      10'd313: inv_x_count_prev = 16'b0000000011010001; // 1/313 = 0.0031948882
      10'd314: inv_x_count_prev = 16'b0000000011010001; // 1/314 = 0.0031847134
      10'd315: inv_x_count_prev = 16'b0000000011010000; // 1/315 = 0.0031746032
      10'd316: inv_x_count_prev = 16'b0000000011001111; // 1/316 = 0.0031645570
      10'd317: inv_x_count_prev = 16'b0000000011001111; // 1/317 = 0.0031545741
      10'd318: inv_x_count_prev = 16'b0000000011001110; // 1/318 = 0.0031446541
      10'd319: inv_x_count_prev = 16'b0000000011001101; // 1/319 = 0.0031347962
      10'd320: inv_x_count_prev = 16'b0000000011001101; // 1/320 = 0.0031250000
      10'd321: inv_x_count_prev = 16'b0000000011001100; // 1/321 = 0.0031152648
      10'd322: inv_x_count_prev = 16'b0000000011001100; // 1/322 = 0.0031055901
      10'd323: inv_x_count_prev = 16'b0000000011001011; // 1/323 = 0.0030959752
      10'd324: inv_x_count_prev = 16'b0000000011001010; // 1/324 = 0.0030864198
      10'd325: inv_x_count_prev = 16'b0000000011001010; // 1/325 = 0.0030769231
      10'd326: inv_x_count_prev = 16'b0000000011001001; // 1/326 = 0.0030674847
      10'd327: inv_x_count_prev = 16'b0000000011001000; // 1/327 = 0.0030581040
      10'd328: inv_x_count_prev = 16'b0000000011001000; // 1/328 = 0.0030487805
      10'd329: inv_x_count_prev = 16'b0000000011000111; // 1/329 = 0.0030395137
      10'd330: inv_x_count_prev = 16'b0000000011000111; // 1/330 = 0.0030303030
      10'd331: inv_x_count_prev = 16'b0000000011000110; // 1/331 = 0.0030211480
      10'd332: inv_x_count_prev = 16'b0000000011000101; // 1/332 = 0.0030120482
      10'd333: inv_x_count_prev = 16'b0000000011000101; // 1/333 = 0.0030030030
      10'd334: inv_x_count_prev = 16'b0000000011000100; // 1/334 = 0.0029940120
      10'd335: inv_x_count_prev = 16'b0000000011000100; // 1/335 = 0.0029850746
      10'd336: inv_x_count_prev = 16'b0000000011000011; // 1/336 = 0.0029761905
      10'd337: inv_x_count_prev = 16'b0000000011000010; // 1/337 = 0.0029673591
      10'd338: inv_x_count_prev = 16'b0000000011000010; // 1/338 = 0.0029585799
      10'd339: inv_x_count_prev = 16'b0000000011000001; // 1/339 = 0.0029498525
      10'd340: inv_x_count_prev = 16'b0000000011000001; // 1/340 = 0.0029411765
      10'd341: inv_x_count_prev = 16'b0000000011000000; // 1/341 = 0.0029325513
      10'd342: inv_x_count_prev = 16'b0000000011000000; // 1/342 = 0.0029239766
      10'd343: inv_x_count_prev = 16'b0000000010111111; // 1/343 = 0.0029154519
      10'd344: inv_x_count_prev = 16'b0000000010111111; // 1/344 = 0.0029069767
      10'd345: inv_x_count_prev = 16'b0000000010111110; // 1/345 = 0.0028985507
      10'd346: inv_x_count_prev = 16'b0000000010111101; // 1/346 = 0.0028901734
      10'd347: inv_x_count_prev = 16'b0000000010111101; // 1/347 = 0.0028818444
      10'd348: inv_x_count_prev = 16'b0000000010111100; // 1/348 = 0.0028735632
      10'd349: inv_x_count_prev = 16'b0000000010111100; // 1/349 = 0.0028653295
      10'd350: inv_x_count_prev = 16'b0000000010111011; // 1/350 = 0.0028571429
      10'd351: inv_x_count_prev = 16'b0000000010111011; // 1/351 = 0.0028490028
      10'd352: inv_x_count_prev = 16'b0000000010111010; // 1/352 = 0.0028409091
      10'd353: inv_x_count_prev = 16'b0000000010111010; // 1/353 = 0.0028328612
      10'd354: inv_x_count_prev = 16'b0000000010111001; // 1/354 = 0.0028248588
      10'd355: inv_x_count_prev = 16'b0000000010111001; // 1/355 = 0.0028169014
      10'd356: inv_x_count_prev = 16'b0000000010111000; // 1/356 = 0.0028089888
      10'd357: inv_x_count_prev = 16'b0000000010111000; // 1/357 = 0.0028011204
      10'd358: inv_x_count_prev = 16'b0000000010110111; // 1/358 = 0.0027932961
      10'd359: inv_x_count_prev = 16'b0000000010110111; // 1/359 = 0.0027855153
      10'd360: inv_x_count_prev = 16'b0000000010110110; // 1/360 = 0.0027777778
      10'd361: inv_x_count_prev = 16'b0000000010110110; // 1/361 = 0.0027700831
      10'd362: inv_x_count_prev = 16'b0000000010110101; // 1/362 = 0.0027624309
      10'd363: inv_x_count_prev = 16'b0000000010110101; // 1/363 = 0.0027548209
      10'd364: inv_x_count_prev = 16'b0000000010110100; // 1/364 = 0.0027472527
      10'd365: inv_x_count_prev = 16'b0000000010110100; // 1/365 = 0.0027397260
      10'd366: inv_x_count_prev = 16'b0000000010110011; // 1/366 = 0.0027322404
      10'd367: inv_x_count_prev = 16'b0000000010110011; // 1/367 = 0.0027247956
      10'd368: inv_x_count_prev = 16'b0000000010110010; // 1/368 = 0.0027173913
      10'd369: inv_x_count_prev = 16'b0000000010110010; // 1/369 = 0.0027100271
      10'd370: inv_x_count_prev = 16'b0000000010110001; // 1/370 = 0.0027027027
      10'd371: inv_x_count_prev = 16'b0000000010110001; // 1/371 = 0.0026954178
      10'd372: inv_x_count_prev = 16'b0000000010110000; // 1/372 = 0.0026881720
      10'd373: inv_x_count_prev = 16'b0000000010110000; // 1/373 = 0.0026809651
      10'd374: inv_x_count_prev = 16'b0000000010101111; // 1/374 = 0.0026737968
      10'd375: inv_x_count_prev = 16'b0000000010101111; // 1/375 = 0.0026666667
      10'd376: inv_x_count_prev = 16'b0000000010101110; // 1/376 = 0.0026595745
      10'd377: inv_x_count_prev = 16'b0000000010101110; // 1/377 = 0.0026525199
      10'd378: inv_x_count_prev = 16'b0000000010101101; // 1/378 = 0.0026455026
      10'd379: inv_x_count_prev = 16'b0000000010101101; // 1/379 = 0.0026385224
      10'd380: inv_x_count_prev = 16'b0000000010101100; // 1/380 = 0.0026315789
      10'd381: inv_x_count_prev = 16'b0000000010101100; // 1/381 = 0.0026246719
      10'd382: inv_x_count_prev = 16'b0000000010101100; // 1/382 = 0.0026178010
      10'd383: inv_x_count_prev = 16'b0000000010101011; // 1/383 = 0.0026109661
      10'd384: inv_x_count_prev = 16'b0000000010101011; // 1/384 = 0.0026041667
      10'd385: inv_x_count_prev = 16'b0000000010101010; // 1/385 = 0.0025974026
      10'd386: inv_x_count_prev = 16'b0000000010101010; // 1/386 = 0.0025906736
      10'd387: inv_x_count_prev = 16'b0000000010101001; // 1/387 = 0.0025839793
      10'd388: inv_x_count_prev = 16'b0000000010101001; // 1/388 = 0.0025773196
      10'd389: inv_x_count_prev = 16'b0000000010101000; // 1/389 = 0.0025706941
      10'd390: inv_x_count_prev = 16'b0000000010101000; // 1/390 = 0.0025641026
      10'd391: inv_x_count_prev = 16'b0000000010101000; // 1/391 = 0.0025575448
      10'd392: inv_x_count_prev = 16'b0000000010100111; // 1/392 = 0.0025510204
      10'd393: inv_x_count_prev = 16'b0000000010100111; // 1/393 = 0.0025445293
      10'd394: inv_x_count_prev = 16'b0000000010100110; // 1/394 = 0.0025380711
      10'd395: inv_x_count_prev = 16'b0000000010100110; // 1/395 = 0.0025316456
      10'd396: inv_x_count_prev = 16'b0000000010100101; // 1/396 = 0.0025252525
      10'd397: inv_x_count_prev = 16'b0000000010100101; // 1/397 = 0.0025188917
      10'd398: inv_x_count_prev = 16'b0000000010100101; // 1/398 = 0.0025125628
      10'd399: inv_x_count_prev = 16'b0000000010100100; // 1/399 = 0.0025062657
      10'd400: inv_x_count_prev = 16'b0000000010100100; // 1/400 = 0.0025000000
      10'd401: inv_x_count_prev = 16'b0000000010100011; // 1/401 = 0.0024937656
      10'd402: inv_x_count_prev = 16'b0000000010100011; // 1/402 = 0.0024875622
      10'd403: inv_x_count_prev = 16'b0000000010100011; // 1/403 = 0.0024813896
      10'd404: inv_x_count_prev = 16'b0000000010100010; // 1/404 = 0.0024752475
      10'd405: inv_x_count_prev = 16'b0000000010100010; // 1/405 = 0.0024691358
      10'd406: inv_x_count_prev = 16'b0000000010100001; // 1/406 = 0.0024630542
      10'd407: inv_x_count_prev = 16'b0000000010100001; // 1/407 = 0.0024570025
      10'd408: inv_x_count_prev = 16'b0000000010100001; // 1/408 = 0.0024509804
      10'd409: inv_x_count_prev = 16'b0000000010100000; // 1/409 = 0.0024449878
      10'd410: inv_x_count_prev = 16'b0000000010100000; // 1/410 = 0.0024390244
      10'd411: inv_x_count_prev = 16'b0000000010011111; // 1/411 = 0.0024330900
      10'd412: inv_x_count_prev = 16'b0000000010011111; // 1/412 = 0.0024271845
      10'd413: inv_x_count_prev = 16'b0000000010011111; // 1/413 = 0.0024213075
      10'd414: inv_x_count_prev = 16'b0000000010011110; // 1/414 = 0.0024154589
      10'd415: inv_x_count_prev = 16'b0000000010011110; // 1/415 = 0.0024096386
      10'd416: inv_x_count_prev = 16'b0000000010011110; // 1/416 = 0.0024038462
      10'd417: inv_x_count_prev = 16'b0000000010011101; // 1/417 = 0.0023980815
      10'd418: inv_x_count_prev = 16'b0000000010011101; // 1/418 = 0.0023923445
      10'd419: inv_x_count_prev = 16'b0000000010011100; // 1/419 = 0.0023866348
      10'd420: inv_x_count_prev = 16'b0000000010011100; // 1/420 = 0.0023809524
      10'd421: inv_x_count_prev = 16'b0000000010011100; // 1/421 = 0.0023752969
      10'd422: inv_x_count_prev = 16'b0000000010011011; // 1/422 = 0.0023696682
      10'd423: inv_x_count_prev = 16'b0000000010011011; // 1/423 = 0.0023640662
      10'd424: inv_x_count_prev = 16'b0000000010011011; // 1/424 = 0.0023584906
      10'd425: inv_x_count_prev = 16'b0000000010011010; // 1/425 = 0.0023529412
      10'd426: inv_x_count_prev = 16'b0000000010011010; // 1/426 = 0.0023474178
      10'd427: inv_x_count_prev = 16'b0000000010011001; // 1/427 = 0.0023419204
      10'd428: inv_x_count_prev = 16'b0000000010011001; // 1/428 = 0.0023364486
      10'd429: inv_x_count_prev = 16'b0000000010011001; // 1/429 = 0.0023310023
      10'd430: inv_x_count_prev = 16'b0000000010011000; // 1/430 = 0.0023255814
      10'd431: inv_x_count_prev = 16'b0000000010011000; // 1/431 = 0.0023201856
      10'd432: inv_x_count_prev = 16'b0000000010011000; // 1/432 = 0.0023148148
      10'd433: inv_x_count_prev = 16'b0000000010010111; // 1/433 = 0.0023094688
      10'd434: inv_x_count_prev = 16'b0000000010010111; // 1/434 = 0.0023041475
      10'd435: inv_x_count_prev = 16'b0000000010010111; // 1/435 = 0.0022988506
      10'd436: inv_x_count_prev = 16'b0000000010010110; // 1/436 = 0.0022935780
      10'd437: inv_x_count_prev = 16'b0000000010010110; // 1/437 = 0.0022883295
      10'd438: inv_x_count_prev = 16'b0000000010010110; // 1/438 = 0.0022831050
      10'd439: inv_x_count_prev = 16'b0000000010010101; // 1/439 = 0.0022779043
      10'd440: inv_x_count_prev = 16'b0000000010010101; // 1/440 = 0.0022727273
      10'd441: inv_x_count_prev = 16'b0000000010010101; // 1/441 = 0.0022675737
      10'd442: inv_x_count_prev = 16'b0000000010010100; // 1/442 = 0.0022624434
      10'd443: inv_x_count_prev = 16'b0000000010010100; // 1/443 = 0.0022573363
      10'd444: inv_x_count_prev = 16'b0000000010010100; // 1/444 = 0.0022522523
      10'd445: inv_x_count_prev = 16'b0000000010010011; // 1/445 = 0.0022471910
      10'd446: inv_x_count_prev = 16'b0000000010010011; // 1/446 = 0.0022421525
      10'd447: inv_x_count_prev = 16'b0000000010010011; // 1/447 = 0.0022371365
      10'd448: inv_x_count_prev = 16'b0000000010010010; // 1/448 = 0.0022321429
      10'd449: inv_x_count_prev = 16'b0000000010010010; // 1/449 = 0.0022271715
      10'd450: inv_x_count_prev = 16'b0000000010010010; // 1/450 = 0.0022222222
      10'd451: inv_x_count_prev = 16'b0000000010010001; // 1/451 = 0.0022172949
      10'd452: inv_x_count_prev = 16'b0000000010010001; // 1/452 = 0.0022123894
      10'd453: inv_x_count_prev = 16'b0000000010010001; // 1/453 = 0.0022075055
      10'd454: inv_x_count_prev = 16'b0000000010010000; // 1/454 = 0.0022026432
      10'd455: inv_x_count_prev = 16'b0000000010010000; // 1/455 = 0.0021978022
      10'd456: inv_x_count_prev = 16'b0000000010010000; // 1/456 = 0.0021929825
      10'd457: inv_x_count_prev = 16'b0000000010001111; // 1/457 = 0.0021881838
      10'd458: inv_x_count_prev = 16'b0000000010001111; // 1/458 = 0.0021834061
      10'd459: inv_x_count_prev = 16'b0000000010001111; // 1/459 = 0.0021786492
      10'd460: inv_x_count_prev = 16'b0000000010001110; // 1/460 = 0.0021739130
      10'd461: inv_x_count_prev = 16'b0000000010001110; // 1/461 = 0.0021691974
      10'd462: inv_x_count_prev = 16'b0000000010001110; // 1/462 = 0.0021645022
      10'd463: inv_x_count_prev = 16'b0000000010001110; // 1/463 = 0.0021598272
      10'd464: inv_x_count_prev = 16'b0000000010001101; // 1/464 = 0.0021551724
      10'd465: inv_x_count_prev = 16'b0000000010001101; // 1/465 = 0.0021505376
      10'd466: inv_x_count_prev = 16'b0000000010001101; // 1/466 = 0.0021459227
      10'd467: inv_x_count_prev = 16'b0000000010001100; // 1/467 = 0.0021413276
      10'd468: inv_x_count_prev = 16'b0000000010001100; // 1/468 = 0.0021367521
      10'd469: inv_x_count_prev = 16'b0000000010001100; // 1/469 = 0.0021321962
      10'd470: inv_x_count_prev = 16'b0000000010001011; // 1/470 = 0.0021276596
      10'd471: inv_x_count_prev = 16'b0000000010001011; // 1/471 = 0.0021231423
      10'd472: inv_x_count_prev = 16'b0000000010001011; // 1/472 = 0.0021186441
      10'd473: inv_x_count_prev = 16'b0000000010001011; // 1/473 = 0.0021141649
      10'd474: inv_x_count_prev = 16'b0000000010001010; // 1/474 = 0.0021097046
      10'd475: inv_x_count_prev = 16'b0000000010001010; // 1/475 = 0.0021052632
      10'd476: inv_x_count_prev = 16'b0000000010001010; // 1/476 = 0.0021008403
      10'd477: inv_x_count_prev = 16'b0000000010001001; // 1/477 = 0.0020964361
      10'd478: inv_x_count_prev = 16'b0000000010001001; // 1/478 = 0.0020920502
      10'd479: inv_x_count_prev = 16'b0000000010001001; // 1/479 = 0.0020876827
      10'd480: inv_x_count_prev = 16'b0000000010001001; // 1/480 = 0.0020833333
      10'd481: inv_x_count_prev = 16'b0000000010001000; // 1/481 = 0.0020790021
      10'd482: inv_x_count_prev = 16'b0000000010001000; // 1/482 = 0.0020746888
      10'd483: inv_x_count_prev = 16'b0000000010001000; // 1/483 = 0.0020703934
      10'd484: inv_x_count_prev = 16'b0000000010000111; // 1/484 = 0.0020661157
      10'd485: inv_x_count_prev = 16'b0000000010000111; // 1/485 = 0.0020618557
      10'd486: inv_x_count_prev = 16'b0000000010000111; // 1/486 = 0.0020576132
      10'd487: inv_x_count_prev = 16'b0000000010000111; // 1/487 = 0.0020533881
      10'd488: inv_x_count_prev = 16'b0000000010000110; // 1/488 = 0.0020491803
      10'd489: inv_x_count_prev = 16'b0000000010000110; // 1/489 = 0.0020449898
      10'd490: inv_x_count_prev = 16'b0000000010000110; // 1/490 = 0.0020408163
      10'd491: inv_x_count_prev = 16'b0000000010000101; // 1/491 = 0.0020366599
      10'd492: inv_x_count_prev = 16'b0000000010000101; // 1/492 = 0.0020325203
      10'd493: inv_x_count_prev = 16'b0000000010000101; // 1/493 = 0.0020283976
      10'd494: inv_x_count_prev = 16'b0000000010000101; // 1/494 = 0.0020242915
      10'd495: inv_x_count_prev = 16'b0000000010000100; // 1/495 = 0.0020202020
      10'd496: inv_x_count_prev = 16'b0000000010000100; // 1/496 = 0.0020161290
      10'd497: inv_x_count_prev = 16'b0000000010000100; // 1/497 = 0.0020120724
      10'd498: inv_x_count_prev = 16'b0000000010000100; // 1/498 = 0.0020080321
      10'd499: inv_x_count_prev = 16'b0000000010000011; // 1/499 = 0.0020040080
      10'd500: inv_x_count_prev = 16'b0000000010000011; // 1/500 = 0.0020000000
      10'd501: inv_x_count_prev = 16'b0000000010000011; // 1/501 = 0.0019960080
      10'd502: inv_x_count_prev = 16'b0000000010000011; // 1/502 = 0.0019920319
      10'd503: inv_x_count_prev = 16'b0000000010000010; // 1/503 = 0.0019880716
      10'd504: inv_x_count_prev = 16'b0000000010000010; // 1/504 = 0.0019841270
      10'd505: inv_x_count_prev = 16'b0000000010000010; // 1/505 = 0.0019801980
      10'd506: inv_x_count_prev = 16'b0000000010000010; // 1/506 = 0.0019762846
      10'd507: inv_x_count_prev = 16'b0000000010000001; // 1/507 = 0.0019723866
      10'd508: inv_x_count_prev = 16'b0000000010000001; // 1/508 = 0.0019685039
      10'd509: inv_x_count_prev = 16'b0000000010000001; // 1/509 = 0.0019646365
      10'd510: inv_x_count_prev = 16'b0000000010000001; // 1/510 = 0.0019607843
      10'd511: inv_x_count_prev = 16'b0000000010000000; // 1/511 = 0.0019569472
      10'd512: inv_x_count_prev = 16'b0000000010000000; // 1/512 = 0.0019531250
      10'd513: inv_x_count_prev = 16'b0000000010000000; // 1/513 = 0.0019493177
      10'd514: inv_x_count_prev = 16'b0000000010000000; // 1/514 = 0.0019455253
      10'd515: inv_x_count_prev = 16'b0000000001111111; // 1/515 = 0.0019417476
      10'd516: inv_x_count_prev = 16'b0000000001111111; // 1/516 = 0.0019379845
      10'd517: inv_x_count_prev = 16'b0000000001111111; // 1/517 = 0.0019342360
      10'd518: inv_x_count_prev = 16'b0000000001111111; // 1/518 = 0.0019305019
      10'd519: inv_x_count_prev = 16'b0000000001111110; // 1/519 = 0.0019267823
      10'd520: inv_x_count_prev = 16'b0000000001111110; // 1/520 = 0.0019230769
      10'd521: inv_x_count_prev = 16'b0000000001111110; // 1/521 = 0.0019193858
      10'd522: inv_x_count_prev = 16'b0000000001111110; // 1/522 = 0.0019157088
      10'd523: inv_x_count_prev = 16'b0000000001111101; // 1/523 = 0.0019120459
      10'd524: inv_x_count_prev = 16'b0000000001111101; // 1/524 = 0.0019083969
      10'd525: inv_x_count_prev = 16'b0000000001111101; // 1/525 = 0.0019047619
      10'd526: inv_x_count_prev = 16'b0000000001111101; // 1/526 = 0.0019011407
      10'd527: inv_x_count_prev = 16'b0000000001111100; // 1/527 = 0.0018975332
      10'd528: inv_x_count_prev = 16'b0000000001111100; // 1/528 = 0.0018939394
      10'd529: inv_x_count_prev = 16'b0000000001111100; // 1/529 = 0.0018903592
      10'd530: inv_x_count_prev = 16'b0000000001111100; // 1/530 = 0.0018867925
      10'd531: inv_x_count_prev = 16'b0000000001111011; // 1/531 = 0.0018832392
      10'd532: inv_x_count_prev = 16'b0000000001111011; // 1/532 = 0.0018796992
      10'd533: inv_x_count_prev = 16'b0000000001111011; // 1/533 = 0.0018761726
      10'd534: inv_x_count_prev = 16'b0000000001111011; // 1/534 = 0.0018726592
      10'd535: inv_x_count_prev = 16'b0000000001111010; // 1/535 = 0.0018691589
      10'd536: inv_x_count_prev = 16'b0000000001111010; // 1/536 = 0.0018656716
      10'd537: inv_x_count_prev = 16'b0000000001111010; // 1/537 = 0.0018621974
      10'd538: inv_x_count_prev = 16'b0000000001111010; // 1/538 = 0.0018587361
      10'd539: inv_x_count_prev = 16'b0000000001111010; // 1/539 = 0.0018552876
      10'd540: inv_x_count_prev = 16'b0000000001111001; // 1/540 = 0.0018518519
      10'd541: inv_x_count_prev = 16'b0000000001111001; // 1/541 = 0.0018484288
      10'd542: inv_x_count_prev = 16'b0000000001111001; // 1/542 = 0.0018450185
      10'd543: inv_x_count_prev = 16'b0000000001111001; // 1/543 = 0.0018416206
      10'd544: inv_x_count_prev = 16'b0000000001111000; // 1/544 = 0.0018382353
      10'd545: inv_x_count_prev = 16'b0000000001111000; // 1/545 = 0.0018348624
      10'd546: inv_x_count_prev = 16'b0000000001111000; // 1/546 = 0.0018315018
      10'd547: inv_x_count_prev = 16'b0000000001111000; // 1/547 = 0.0018281536
      10'd548: inv_x_count_prev = 16'b0000000001111000; // 1/548 = 0.0018248175
      10'd549: inv_x_count_prev = 16'b0000000001110111; // 1/549 = 0.0018214936
      10'd550: inv_x_count_prev = 16'b0000000001110111; // 1/550 = 0.0018181818
      10'd551: inv_x_count_prev = 16'b0000000001110111; // 1/551 = 0.0018148820
      10'd552: inv_x_count_prev = 16'b0000000001110111; // 1/552 = 0.0018115942
      10'd553: inv_x_count_prev = 16'b0000000001110111; // 1/553 = 0.0018083183
      10'd554: inv_x_count_prev = 16'b0000000001110110; // 1/554 = 0.0018050542
      10'd555: inv_x_count_prev = 16'b0000000001110110; // 1/555 = 0.0018018018
      10'd556: inv_x_count_prev = 16'b0000000001110110; // 1/556 = 0.0017985612
      10'd557: inv_x_count_prev = 16'b0000000001110110; // 1/557 = 0.0017953321
      10'd558: inv_x_count_prev = 16'b0000000001110101; // 1/558 = 0.0017921147
      10'd559: inv_x_count_prev = 16'b0000000001110101; // 1/559 = 0.0017889088
      10'd560: inv_x_count_prev = 16'b0000000001110101; // 1/560 = 0.0017857143
      10'd561: inv_x_count_prev = 16'b0000000001110101; // 1/561 = 0.0017825312
      10'd562: inv_x_count_prev = 16'b0000000001110101; // 1/562 = 0.0017793594
      10'd563: inv_x_count_prev = 16'b0000000001110100; // 1/563 = 0.0017761989
      10'd564: inv_x_count_prev = 16'b0000000001110100; // 1/564 = 0.0017730496
      10'd565: inv_x_count_prev = 16'b0000000001110100; // 1/565 = 0.0017699115
      10'd566: inv_x_count_prev = 16'b0000000001110100; // 1/566 = 0.0017667845
      10'd567: inv_x_count_prev = 16'b0000000001110100; // 1/567 = 0.0017636684
      10'd568: inv_x_count_prev = 16'b0000000001110011; // 1/568 = 0.0017605634
      10'd569: inv_x_count_prev = 16'b0000000001110011; // 1/569 = 0.0017574692
      10'd570: inv_x_count_prev = 16'b0000000001110011; // 1/570 = 0.0017543860
      10'd571: inv_x_count_prev = 16'b0000000001110011; // 1/571 = 0.0017513135
      10'd572: inv_x_count_prev = 16'b0000000001110011; // 1/572 = 0.0017482517
      10'd573: inv_x_count_prev = 16'b0000000001110010; // 1/573 = 0.0017452007
      10'd574: inv_x_count_prev = 16'b0000000001110010; // 1/574 = 0.0017421603
      10'd575: inv_x_count_prev = 16'b0000000001110010; // 1/575 = 0.0017391304
      10'd576: inv_x_count_prev = 16'b0000000001110010; // 1/576 = 0.0017361111
      10'd577: inv_x_count_prev = 16'b0000000001110010; // 1/577 = 0.0017331023
      10'd578: inv_x_count_prev = 16'b0000000001110001; // 1/578 = 0.0017301038
      10'd579: inv_x_count_prev = 16'b0000000001110001; // 1/579 = 0.0017271157
      10'd580: inv_x_count_prev = 16'b0000000001110001; // 1/580 = 0.0017241379
      10'd581: inv_x_count_prev = 16'b0000000001110001; // 1/581 = 0.0017211704
      10'd582: inv_x_count_prev = 16'b0000000001110001; // 1/582 = 0.0017182131
      10'd583: inv_x_count_prev = 16'b0000000001110000; // 1/583 = 0.0017152659
      10'd584: inv_x_count_prev = 16'b0000000001110000; // 1/584 = 0.0017123288
      10'd585: inv_x_count_prev = 16'b0000000001110000; // 1/585 = 0.0017094017
      10'd586: inv_x_count_prev = 16'b0000000001110000; // 1/586 = 0.0017064846
      10'd587: inv_x_count_prev = 16'b0000000001110000; // 1/587 = 0.0017035775
      10'd588: inv_x_count_prev = 16'b0000000001101111; // 1/588 = 0.0017006803
      10'd589: inv_x_count_prev = 16'b0000000001101111; // 1/589 = 0.0016977929
      10'd590: inv_x_count_prev = 16'b0000000001101111; // 1/590 = 0.0016949153
      10'd591: inv_x_count_prev = 16'b0000000001101111; // 1/591 = 0.0016920474
      10'd592: inv_x_count_prev = 16'b0000000001101111; // 1/592 = 0.0016891892
      10'd593: inv_x_count_prev = 16'b0000000001101111; // 1/593 = 0.0016863406
      10'd594: inv_x_count_prev = 16'b0000000001101110; // 1/594 = 0.0016835017
      10'd595: inv_x_count_prev = 16'b0000000001101110; // 1/595 = 0.0016806723
      10'd596: inv_x_count_prev = 16'b0000000001101110; // 1/596 = 0.0016778523
      10'd597: inv_x_count_prev = 16'b0000000001101110; // 1/597 = 0.0016750419
      10'd598: inv_x_count_prev = 16'b0000000001101110; // 1/598 = 0.0016722408
      10'd599: inv_x_count_prev = 16'b0000000001101101; // 1/599 = 0.0016694491
      10'd600: inv_x_count_prev = 16'b0000000001101101; // 1/600 = 0.0016666667
      10'd601: inv_x_count_prev = 16'b0000000001101101; // 1/601 = 0.0016638935
      10'd602: inv_x_count_prev = 16'b0000000001101101; // 1/602 = 0.0016611296
      10'd603: inv_x_count_prev = 16'b0000000001101101; // 1/603 = 0.0016583748
      10'd604: inv_x_count_prev = 16'b0000000001101101; // 1/604 = 0.0016556291
      10'd605: inv_x_count_prev = 16'b0000000001101100; // 1/605 = 0.0016528926
      10'd606: inv_x_count_prev = 16'b0000000001101100; // 1/606 = 0.0016501650
      10'd607: inv_x_count_prev = 16'b0000000001101100; // 1/607 = 0.0016474465
      10'd608: inv_x_count_prev = 16'b0000000001101100; // 1/608 = 0.0016447368
      10'd609: inv_x_count_prev = 16'b0000000001101100; // 1/609 = 0.0016420361
      10'd610: inv_x_count_prev = 16'b0000000001101011; // 1/610 = 0.0016393443
      10'd611: inv_x_count_prev = 16'b0000000001101011; // 1/611 = 0.0016366612
      10'd612: inv_x_count_prev = 16'b0000000001101011; // 1/612 = 0.0016339869
      10'd613: inv_x_count_prev = 16'b0000000001101011; // 1/613 = 0.0016313214
      10'd614: inv_x_count_prev = 16'b0000000001101011; // 1/614 = 0.0016286645
      10'd615: inv_x_count_prev = 16'b0000000001101011; // 1/615 = 0.0016260163
      10'd616: inv_x_count_prev = 16'b0000000001101010; // 1/616 = 0.0016233766
      10'd617: inv_x_count_prev = 16'b0000000001101010; // 1/617 = 0.0016207455
      10'd618: inv_x_count_prev = 16'b0000000001101010; // 1/618 = 0.0016181230
      10'd619: inv_x_count_prev = 16'b0000000001101010; // 1/619 = 0.0016155089
      10'd620: inv_x_count_prev = 16'b0000000001101010; // 1/620 = 0.0016129032
      10'd621: inv_x_count_prev = 16'b0000000001101010; // 1/621 = 0.0016103060
      10'd622: inv_x_count_prev = 16'b0000000001101001; // 1/622 = 0.0016077170
      10'd623: inv_x_count_prev = 16'b0000000001101001; // 1/623 = 0.0016051364
      10'd624: inv_x_count_prev = 16'b0000000001101001; // 1/624 = 0.0016025641
      10'd625: inv_x_count_prev = 16'b0000000001101001; // 1/625 = 0.0016000000
      10'd626: inv_x_count_prev = 16'b0000000001101001; // 1/626 = 0.0015974441
      10'd627: inv_x_count_prev = 16'b0000000001101001; // 1/627 = 0.0015948963
      10'd628: inv_x_count_prev = 16'b0000000001101000; // 1/628 = 0.0015923567
      10'd629: inv_x_count_prev = 16'b0000000001101000; // 1/629 = 0.0015898251
      10'd630: inv_x_count_prev = 16'b0000000001101000; // 1/630 = 0.0015873016
      10'd631: inv_x_count_prev = 16'b0000000001101000; // 1/631 = 0.0015847861
      10'd632: inv_x_count_prev = 16'b0000000001101000; // 1/632 = 0.0015822785
      10'd633: inv_x_count_prev = 16'b0000000001101000; // 1/633 = 0.0015797788
      10'd634: inv_x_count_prev = 16'b0000000001100111; // 1/634 = 0.0015772871
      10'd635: inv_x_count_prev = 16'b0000000001100111; // 1/635 = 0.0015748031
      10'd636: inv_x_count_prev = 16'b0000000001100111; // 1/636 = 0.0015723270
      10'd637: inv_x_count_prev = 16'b0000000001100111; // 1/637 = 0.0015698587
      10'd638: inv_x_count_prev = 16'b0000000001100111; // 1/638 = 0.0015673981
      10'd639: inv_x_count_prev = 16'b0000000001100111; // 1/639 = 0.0015649452
      10'd640: inv_x_count_prev = 16'b0000000001100110; // 1/640 = 0.0015625000
      10'd641: inv_x_count_prev = 16'b0000000001100110; // 1/641 = 0.0015600624
      10'd642: inv_x_count_prev = 16'b0000000001100110; // 1/642 = 0.0015576324
      10'd643: inv_x_count_prev = 16'b0000000001100110; // 1/643 = 0.0015552100
      10'd644: inv_x_count_prev = 16'b0000000001100110; // 1/644 = 0.0015527950
      10'd645: inv_x_count_prev = 16'b0000000001100110; // 1/645 = 0.0015503876
      10'd646: inv_x_count_prev = 16'b0000000001100101; // 1/646 = 0.0015479876
      10'd647: inv_x_count_prev = 16'b0000000001100101; // 1/647 = 0.0015455951
      10'd648: inv_x_count_prev = 16'b0000000001100101; // 1/648 = 0.0015432099
      10'd649: inv_x_count_prev = 16'b0000000001100101; // 1/649 = 0.0015408320
      10'd650: inv_x_count_prev = 16'b0000000001100101; // 1/650 = 0.0015384615
      10'd651: inv_x_count_prev = 16'b0000000001100101; // 1/651 = 0.0015360983
      10'd652: inv_x_count_prev = 16'b0000000001100101; // 1/652 = 0.0015337423
      10'd653: inv_x_count_prev = 16'b0000000001100100; // 1/653 = 0.0015313936
      10'd654: inv_x_count_prev = 16'b0000000001100100; // 1/654 = 0.0015290520
      10'd655: inv_x_count_prev = 16'b0000000001100100; // 1/655 = 0.0015267176
      10'd656: inv_x_count_prev = 16'b0000000001100100; // 1/656 = 0.0015243902
      10'd657: inv_x_count_prev = 16'b0000000001100100; // 1/657 = 0.0015220700
      10'd658: inv_x_count_prev = 16'b0000000001100100; // 1/658 = 0.0015197568
      10'd659: inv_x_count_prev = 16'b0000000001100011; // 1/659 = 0.0015174507
      10'd660: inv_x_count_prev = 16'b0000000001100011; // 1/660 = 0.0015151515
      10'd661: inv_x_count_prev = 16'b0000000001100011; // 1/661 = 0.0015128593
      10'd662: inv_x_count_prev = 16'b0000000001100011; // 1/662 = 0.0015105740
      10'd663: inv_x_count_prev = 16'b0000000001100011; // 1/663 = 0.0015082956
      10'd664: inv_x_count_prev = 16'b0000000001100011; // 1/664 = 0.0015060241
      10'd665: inv_x_count_prev = 16'b0000000001100011; // 1/665 = 0.0015037594
      10'd666: inv_x_count_prev = 16'b0000000001100010; // 1/666 = 0.0015015015
      10'd667: inv_x_count_prev = 16'b0000000001100010; // 1/667 = 0.0014992504
      10'd668: inv_x_count_prev = 16'b0000000001100010; // 1/668 = 0.0014970060
      10'd669: inv_x_count_prev = 16'b0000000001100010; // 1/669 = 0.0014947683
      10'd670: inv_x_count_prev = 16'b0000000001100010; // 1/670 = 0.0014925373
      10'd671: inv_x_count_prev = 16'b0000000001100010; // 1/671 = 0.0014903130
      10'd672: inv_x_count_prev = 16'b0000000001100010; // 1/672 = 0.0014880952
      10'd673: inv_x_count_prev = 16'b0000000001100001; // 1/673 = 0.0014858841
      10'd674: inv_x_count_prev = 16'b0000000001100001; // 1/674 = 0.0014836795
      10'd675: inv_x_count_prev = 16'b0000000001100001; // 1/675 = 0.0014814815
      10'd676: inv_x_count_prev = 16'b0000000001100001; // 1/676 = 0.0014792899
      10'd677: inv_x_count_prev = 16'b0000000001100001; // 1/677 = 0.0014771049
      10'd678: inv_x_count_prev = 16'b0000000001100001; // 1/678 = 0.0014749263
      10'd679: inv_x_count_prev = 16'b0000000001100001; // 1/679 = 0.0014727541
      10'd680: inv_x_count_prev = 16'b0000000001100000; // 1/680 = 0.0014705882
      10'd681: inv_x_count_prev = 16'b0000000001100000; // 1/681 = 0.0014684288
      10'd682: inv_x_count_prev = 16'b0000000001100000; // 1/682 = 0.0014662757
      10'd683: inv_x_count_prev = 16'b0000000001100000; // 1/683 = 0.0014641288
      10'd684: inv_x_count_prev = 16'b0000000001100000; // 1/684 = 0.0014619883
      10'd685: inv_x_count_prev = 16'b0000000001100000; // 1/685 = 0.0014598540
      10'd686: inv_x_count_prev = 16'b0000000001100000; // 1/686 = 0.0014577259
      10'd687: inv_x_count_prev = 16'b0000000001011111; // 1/687 = 0.0014556041
      10'd688: inv_x_count_prev = 16'b0000000001011111; // 1/688 = 0.0014534884
      10'd689: inv_x_count_prev = 16'b0000000001011111; // 1/689 = 0.0014513788
      10'd690: inv_x_count_prev = 16'b0000000001011111; // 1/690 = 0.0014492754
      10'd691: inv_x_count_prev = 16'b0000000001011111; // 1/691 = 0.0014471780
      10'd692: inv_x_count_prev = 16'b0000000001011111; // 1/692 = 0.0014450867
      10'd693: inv_x_count_prev = 16'b0000000001011111; // 1/693 = 0.0014430014
      10'd694: inv_x_count_prev = 16'b0000000001011110; // 1/694 = 0.0014409222
      10'd695: inv_x_count_prev = 16'b0000000001011110; // 1/695 = 0.0014388489
      10'd696: inv_x_count_prev = 16'b0000000001011110; // 1/696 = 0.0014367816
      10'd697: inv_x_count_prev = 16'b0000000001011110; // 1/697 = 0.0014347202
      10'd698: inv_x_count_prev = 16'b0000000001011110; // 1/698 = 0.0014326648
      10'd699: inv_x_count_prev = 16'b0000000001011110; // 1/699 = 0.0014306152
      10'd700: inv_x_count_prev = 16'b0000000001011110; // 1/700 = 0.0014285714
      10'd701: inv_x_count_prev = 16'b0000000001011101; // 1/701 = 0.0014265335
      10'd702: inv_x_count_prev = 16'b0000000001011101; // 1/702 = 0.0014245014
      10'd703: inv_x_count_prev = 16'b0000000001011101; // 1/703 = 0.0014224751
      10'd704: inv_x_count_prev = 16'b0000000001011101; // 1/704 = 0.0014204545
      10'd705: inv_x_count_prev = 16'b0000000001011101; // 1/705 = 0.0014184397
      10'd706: inv_x_count_prev = 16'b0000000001011101; // 1/706 = 0.0014164306
      10'd707: inv_x_count_prev = 16'b0000000001011101; // 1/707 = 0.0014144272
      10'd708: inv_x_count_prev = 16'b0000000001011101; // 1/708 = 0.0014124294
      10'd709: inv_x_count_prev = 16'b0000000001011100; // 1/709 = 0.0014104372
      10'd710: inv_x_count_prev = 16'b0000000001011100; // 1/710 = 0.0014084507
      10'd711: inv_x_count_prev = 16'b0000000001011100; // 1/711 = 0.0014064698
      10'd712: inv_x_count_prev = 16'b0000000001011100; // 1/712 = 0.0014044944
      10'd713: inv_x_count_prev = 16'b0000000001011100; // 1/713 = 0.0014025245
      10'd714: inv_x_count_prev = 16'b0000000001011100; // 1/714 = 0.0014005602
      10'd715: inv_x_count_prev = 16'b0000000001011100; // 1/715 = 0.0013986014
      10'd716: inv_x_count_prev = 16'b0000000001011100; // 1/716 = 0.0013966480
      10'd717: inv_x_count_prev = 16'b0000000001011011; // 1/717 = 0.0013947001
      10'd718: inv_x_count_prev = 16'b0000000001011011; // 1/718 = 0.0013927577
      10'd719: inv_x_count_prev = 16'b0000000001011011; // 1/719 = 0.0013908206
      10'd720: inv_x_count_prev = 16'b0000000001011011; // 1/720 = 0.0013888889
      10'd721: inv_x_count_prev = 16'b0000000001011011; // 1/721 = 0.0013869626
      10'd722: inv_x_count_prev = 16'b0000000001011011; // 1/722 = 0.0013850416
      10'd723: inv_x_count_prev = 16'b0000000001011011; // 1/723 = 0.0013831259
      10'd724: inv_x_count_prev = 16'b0000000001011011; // 1/724 = 0.0013812155
      10'd725: inv_x_count_prev = 16'b0000000001011010; // 1/725 = 0.0013793103
      10'd726: inv_x_count_prev = 16'b0000000001011010; // 1/726 = 0.0013774105
      10'd727: inv_x_count_prev = 16'b0000000001011010; // 1/727 = 0.0013755158
      10'd728: inv_x_count_prev = 16'b0000000001011010; // 1/728 = 0.0013736264
      10'd729: inv_x_count_prev = 16'b0000000001011010; // 1/729 = 0.0013717421
      10'd730: inv_x_count_prev = 16'b0000000001011010; // 1/730 = 0.0013698630
      10'd731: inv_x_count_prev = 16'b0000000001011010; // 1/731 = 0.0013679891
      10'd732: inv_x_count_prev = 16'b0000000001011010; // 1/732 = 0.0013661202
      10'd733: inv_x_count_prev = 16'b0000000001011001; // 1/733 = 0.0013642565
      10'd734: inv_x_count_prev = 16'b0000000001011001; // 1/734 = 0.0013623978
      10'd735: inv_x_count_prev = 16'b0000000001011001; // 1/735 = 0.0013605442
      10'd736: inv_x_count_prev = 16'b0000000001011001; // 1/736 = 0.0013586957
      10'd737: inv_x_count_prev = 16'b0000000001011001; // 1/737 = 0.0013568521
      10'd738: inv_x_count_prev = 16'b0000000001011001; // 1/738 = 0.0013550136
      10'd739: inv_x_count_prev = 16'b0000000001011001; // 1/739 = 0.0013531800
      10'd740: inv_x_count_prev = 16'b0000000001011001; // 1/740 = 0.0013513514
      10'd741: inv_x_count_prev = 16'b0000000001011000; // 1/741 = 0.0013495277
      10'd742: inv_x_count_prev = 16'b0000000001011000; // 1/742 = 0.0013477089
      10'd743: inv_x_count_prev = 16'b0000000001011000; // 1/743 = 0.0013458950
      10'd744: inv_x_count_prev = 16'b0000000001011000; // 1/744 = 0.0013440860
      10'd745: inv_x_count_prev = 16'b0000000001011000; // 1/745 = 0.0013422819
      10'd746: inv_x_count_prev = 16'b0000000001011000; // 1/746 = 0.0013404826
      10'd747: inv_x_count_prev = 16'b0000000001011000; // 1/747 = 0.0013386881
      10'd748: inv_x_count_prev = 16'b0000000001011000; // 1/748 = 0.0013368984
      10'd749: inv_x_count_prev = 16'b0000000001010111; // 1/749 = 0.0013351135
      10'd750: inv_x_count_prev = 16'b0000000001010111; // 1/750 = 0.0013333333
      10'd751: inv_x_count_prev = 16'b0000000001010111; // 1/751 = 0.0013315579
      10'd752: inv_x_count_prev = 16'b0000000001010111; // 1/752 = 0.0013297872
      10'd753: inv_x_count_prev = 16'b0000000001010111; // 1/753 = 0.0013280212
      10'd754: inv_x_count_prev = 16'b0000000001010111; // 1/754 = 0.0013262599
      10'd755: inv_x_count_prev = 16'b0000000001010111; // 1/755 = 0.0013245033
      10'd756: inv_x_count_prev = 16'b0000000001010111; // 1/756 = 0.0013227513
      10'd757: inv_x_count_prev = 16'b0000000001010111; // 1/757 = 0.0013210040
      10'd758: inv_x_count_prev = 16'b0000000001010110; // 1/758 = 0.0013192612
      10'd759: inv_x_count_prev = 16'b0000000001010110; // 1/759 = 0.0013175231
      10'd760: inv_x_count_prev = 16'b0000000001010110; // 1/760 = 0.0013157895
      10'd761: inv_x_count_prev = 16'b0000000001010110; // 1/761 = 0.0013140604
      10'd762: inv_x_count_prev = 16'b0000000001010110; // 1/762 = 0.0013123360
      10'd763: inv_x_count_prev = 16'b0000000001010110; // 1/763 = 0.0013106160
      10'd764: inv_x_count_prev = 16'b0000000001010110; // 1/764 = 0.0013089005
      10'd765: inv_x_count_prev = 16'b0000000001010110; // 1/765 = 0.0013071895
      10'd766: inv_x_count_prev = 16'b0000000001010110; // 1/766 = 0.0013054830
      10'd767: inv_x_count_prev = 16'b0000000001010101; // 1/767 = 0.0013037810
      10'd768: inv_x_count_prev = 16'b0000000001010101; // 1/768 = 0.0013020833
      10'd769: inv_x_count_prev = 16'b0000000001010101; // 1/769 = 0.0013003901
      10'd770: inv_x_count_prev = 16'b0000000001010101; // 1/770 = 0.0012987013
      10'd771: inv_x_count_prev = 16'b0000000001010101; // 1/771 = 0.0012970169
      10'd772: inv_x_count_prev = 16'b0000000001010101; // 1/772 = 0.0012953368
      10'd773: inv_x_count_prev = 16'b0000000001010101; // 1/773 = 0.0012936611
      10'd774: inv_x_count_prev = 16'b0000000001010101; // 1/774 = 0.0012919897
      10'd775: inv_x_count_prev = 16'b0000000001010101; // 1/775 = 0.0012903226
      10'd776: inv_x_count_prev = 16'b0000000001010100; // 1/776 = 0.0012886598
      10'd777: inv_x_count_prev = 16'b0000000001010100; // 1/777 = 0.0012870013
      10'd778: inv_x_count_prev = 16'b0000000001010100; // 1/778 = 0.0012853470
      10'd779: inv_x_count_prev = 16'b0000000001010100; // 1/779 = 0.0012836970
      10'd780: inv_x_count_prev = 16'b0000000001010100; // 1/780 = 0.0012820513
      10'd781: inv_x_count_prev = 16'b0000000001010100; // 1/781 = 0.0012804097
      10'd782: inv_x_count_prev = 16'b0000000001010100; // 1/782 = 0.0012787724
      10'd783: inv_x_count_prev = 16'b0000000001010100; // 1/783 = 0.0012771392
      10'd784: inv_x_count_prev = 16'b0000000001010100; // 1/784 = 0.0012755102
      10'd785: inv_x_count_prev = 16'b0000000001010011; // 1/785 = 0.0012738854
      10'd786: inv_x_count_prev = 16'b0000000001010011; // 1/786 = 0.0012722646
      10'd787: inv_x_count_prev = 16'b0000000001010011; // 1/787 = 0.0012706480
      10'd788: inv_x_count_prev = 16'b0000000001010011; // 1/788 = 0.0012690355
      10'd789: inv_x_count_prev = 16'b0000000001010011; // 1/789 = 0.0012674271
      10'd790: inv_x_count_prev = 16'b0000000001010011; // 1/790 = 0.0012658228
      10'd791: inv_x_count_prev = 16'b0000000001010011; // 1/791 = 0.0012642225
      10'd792: inv_x_count_prev = 16'b0000000001010011; // 1/792 = 0.0012626263
      10'd793: inv_x_count_prev = 16'b0000000001010011; // 1/793 = 0.0012610340
      10'd794: inv_x_count_prev = 16'b0000000001010011; // 1/794 = 0.0012594458
      10'd795: inv_x_count_prev = 16'b0000000001010010; // 1/795 = 0.0012578616
      10'd796: inv_x_count_prev = 16'b0000000001010010; // 1/796 = 0.0012562814
      10'd797: inv_x_count_prev = 16'b0000000001010010; // 1/797 = 0.0012547051
      10'd798: inv_x_count_prev = 16'b0000000001010010; // 1/798 = 0.0012531328
      10'd799: inv_x_count_prev = 16'b0000000001010010; // 1/799 = 0.0012515645
      10'd800: inv_x_count_prev = 16'b0000000001010010; // 1/800 = 0.0012500000
      10'd801: inv_x_count_prev = 16'b0000000001010010; // 1/801 = 0.0012484395
      10'd802: inv_x_count_prev = 16'b0000000001010010; // 1/802 = 0.0012468828
      10'd803: inv_x_count_prev = 16'b0000000001010010; // 1/803 = 0.0012453300
      10'd804: inv_x_count_prev = 16'b0000000001010010; // 1/804 = 0.0012437811
      10'd805: inv_x_count_prev = 16'b0000000001010001; // 1/805 = 0.0012422360
      10'd806: inv_x_count_prev = 16'b0000000001010001; // 1/806 = 0.0012406948
      10'd807: inv_x_count_prev = 16'b0000000001010001; // 1/807 = 0.0012391574
      10'd808: inv_x_count_prev = 16'b0000000001010001; // 1/808 = 0.0012376238
      10'd809: inv_x_count_prev = 16'b0000000001010001; // 1/809 = 0.0012360939
      10'd810: inv_x_count_prev = 16'b0000000001010001; // 1/810 = 0.0012345679
      10'd811: inv_x_count_prev = 16'b0000000001010001; // 1/811 = 0.0012330456
      10'd812: inv_x_count_prev = 16'b0000000001010001; // 1/812 = 0.0012315271
      10'd813: inv_x_count_prev = 16'b0000000001010001; // 1/813 = 0.0012300123
      10'd814: inv_x_count_prev = 16'b0000000001010001; // 1/814 = 0.0012285012
      10'd815: inv_x_count_prev = 16'b0000000001010000; // 1/815 = 0.0012269939
      10'd816: inv_x_count_prev = 16'b0000000001010000; // 1/816 = 0.0012254902
      10'd817: inv_x_count_prev = 16'b0000000001010000; // 1/817 = 0.0012239902
      10'd818: inv_x_count_prev = 16'b0000000001010000; // 1/818 = 0.0012224939
      10'd819: inv_x_count_prev = 16'b0000000001010000; // 1/819 = 0.0012210012
      10'd820: inv_x_count_prev = 16'b0000000001010000; // 1/820 = 0.0012195122
      10'd821: inv_x_count_prev = 16'b0000000001010000; // 1/821 = 0.0012180268
      10'd822: inv_x_count_prev = 16'b0000000001010000; // 1/822 = 0.0012165450
      10'd823: inv_x_count_prev = 16'b0000000001010000; // 1/823 = 0.0012150668
      10'd824: inv_x_count_prev = 16'b0000000001010000; // 1/824 = 0.0012135922
      10'd825: inv_x_count_prev = 16'b0000000001001111; // 1/825 = 0.0012121212
      10'd826: inv_x_count_prev = 16'b0000000001001111; // 1/826 = 0.0012106538
      10'd827: inv_x_count_prev = 16'b0000000001001111; // 1/827 = 0.0012091898
      10'd828: inv_x_count_prev = 16'b0000000001001111; // 1/828 = 0.0012077295
      10'd829: inv_x_count_prev = 16'b0000000001001111; // 1/829 = 0.0012062726
      10'd830: inv_x_count_prev = 16'b0000000001001111; // 1/830 = 0.0012048193
      10'd831: inv_x_count_prev = 16'b0000000001001111; // 1/831 = 0.0012033694
      10'd832: inv_x_count_prev = 16'b0000000001001111; // 1/832 = 0.0012019231
      10'd833: inv_x_count_prev = 16'b0000000001001111; // 1/833 = 0.0012004802
      10'd834: inv_x_count_prev = 16'b0000000001001111; // 1/834 = 0.0011990408
      10'd835: inv_x_count_prev = 16'b0000000001001110; // 1/835 = 0.0011976048
      10'd836: inv_x_count_prev = 16'b0000000001001110; // 1/836 = 0.0011961722
      10'd837: inv_x_count_prev = 16'b0000000001001110; // 1/837 = 0.0011947431
      10'd838: inv_x_count_prev = 16'b0000000001001110; // 1/838 = 0.0011933174
      10'd839: inv_x_count_prev = 16'b0000000001001110; // 1/839 = 0.0011918951
      10'd840: inv_x_count_prev = 16'b0000000001001110; // 1/840 = 0.0011904762
      10'd841: inv_x_count_prev = 16'b0000000001001110; // 1/841 = 0.0011890606
      10'd842: inv_x_count_prev = 16'b0000000001001110; // 1/842 = 0.0011876485
      10'd843: inv_x_count_prev = 16'b0000000001001110; // 1/843 = 0.0011862396
      10'd844: inv_x_count_prev = 16'b0000000001001110; // 1/844 = 0.0011848341
      10'd845: inv_x_count_prev = 16'b0000000001001110; // 1/845 = 0.0011834320
      10'd846: inv_x_count_prev = 16'b0000000001001101; // 1/846 = 0.0011820331
      10'd847: inv_x_count_prev = 16'b0000000001001101; // 1/847 = 0.0011806375
      10'd848: inv_x_count_prev = 16'b0000000001001101; // 1/848 = 0.0011792453
      10'd849: inv_x_count_prev = 16'b0000000001001101; // 1/849 = 0.0011778563
      10'd850: inv_x_count_prev = 16'b0000000001001101; // 1/850 = 0.0011764706
      10'd851: inv_x_count_prev = 16'b0000000001001101; // 1/851 = 0.0011750881
      10'd852: inv_x_count_prev = 16'b0000000001001101; // 1/852 = 0.0011737089
      10'd853: inv_x_count_prev = 16'b0000000001001101; // 1/853 = 0.0011723329
      10'd854: inv_x_count_prev = 16'b0000000001001101; // 1/854 = 0.0011709602
      10'd855: inv_x_count_prev = 16'b0000000001001101; // 1/855 = 0.0011695906
      10'd856: inv_x_count_prev = 16'b0000000001001101; // 1/856 = 0.0011682243
      10'd857: inv_x_count_prev = 16'b0000000001001100; // 1/857 = 0.0011668611
      10'd858: inv_x_count_prev = 16'b0000000001001100; // 1/858 = 0.0011655012
      10'd859: inv_x_count_prev = 16'b0000000001001100; // 1/859 = 0.0011641444
      10'd860: inv_x_count_prev = 16'b0000000001001100; // 1/860 = 0.0011627907
      10'd861: inv_x_count_prev = 16'b0000000001001100; // 1/861 = 0.0011614402
      10'd862: inv_x_count_prev = 16'b0000000001001100; // 1/862 = 0.0011600928
      10'd863: inv_x_count_prev = 16'b0000000001001100; // 1/863 = 0.0011587486
      10'd864: inv_x_count_prev = 16'b0000000001001100; // 1/864 = 0.0011574074
      10'd865: inv_x_count_prev = 16'b0000000001001100; // 1/865 = 0.0011560694
      10'd866: inv_x_count_prev = 16'b0000000001001100; // 1/866 = 0.0011547344
      10'd867: inv_x_count_prev = 16'b0000000001001100; // 1/867 = 0.0011534025
      10'd868: inv_x_count_prev = 16'b0000000001001100; // 1/868 = 0.0011520737
      10'd869: inv_x_count_prev = 16'b0000000001001011; // 1/869 = 0.0011507480
      10'd870: inv_x_count_prev = 16'b0000000001001011; // 1/870 = 0.0011494253
      10'd871: inv_x_count_prev = 16'b0000000001001011; // 1/871 = 0.0011481056
      10'd872: inv_x_count_prev = 16'b0000000001001011; // 1/872 = 0.0011467890
      10'd873: inv_x_count_prev = 16'b0000000001001011; // 1/873 = 0.0011454754
      10'd874: inv_x_count_prev = 16'b0000000001001011; // 1/874 = 0.0011441648
      10'd875: inv_x_count_prev = 16'b0000000001001011; // 1/875 = 0.0011428571
      10'd876: inv_x_count_prev = 16'b0000000001001011; // 1/876 = 0.0011415525
      10'd877: inv_x_count_prev = 16'b0000000001001011; // 1/877 = 0.0011402509
      10'd878: inv_x_count_prev = 16'b0000000001001011; // 1/878 = 0.0011389522
      10'd879: inv_x_count_prev = 16'b0000000001001011; // 1/879 = 0.0011376564
      10'd880: inv_x_count_prev = 16'b0000000001001010; // 1/880 = 0.0011363636
      10'd881: inv_x_count_prev = 16'b0000000001001010; // 1/881 = 0.0011350738
      10'd882: inv_x_count_prev = 16'b0000000001001010; // 1/882 = 0.0011337868
      10'd883: inv_x_count_prev = 16'b0000000001001010; // 1/883 = 0.0011325028
      10'd884: inv_x_count_prev = 16'b0000000001001010; // 1/884 = 0.0011312217
      10'd885: inv_x_count_prev = 16'b0000000001001010; // 1/885 = 0.0011299435
      10'd886: inv_x_count_prev = 16'b0000000001001010; // 1/886 = 0.0011286682
      10'd887: inv_x_count_prev = 16'b0000000001001010; // 1/887 = 0.0011273957
      10'd888: inv_x_count_prev = 16'b0000000001001010; // 1/888 = 0.0011261261
      10'd889: inv_x_count_prev = 16'b0000000001001010; // 1/889 = 0.0011248594
      10'd890: inv_x_count_prev = 16'b0000000001001010; // 1/890 = 0.0011235955
      10'd891: inv_x_count_prev = 16'b0000000001001010; // 1/891 = 0.0011223345
      10'd892: inv_x_count_prev = 16'b0000000001001001; // 1/892 = 0.0011210762
      10'd893: inv_x_count_prev = 16'b0000000001001001; // 1/893 = 0.0011198208
      10'd894: inv_x_count_prev = 16'b0000000001001001; // 1/894 = 0.0011185682
      10'd895: inv_x_count_prev = 16'b0000000001001001; // 1/895 = 0.0011173184
      10'd896: inv_x_count_prev = 16'b0000000001001001; // 1/896 = 0.0011160714
      10'd897: inv_x_count_prev = 16'b0000000001001001; // 1/897 = 0.0011148272
      10'd898: inv_x_count_prev = 16'b0000000001001001; // 1/898 = 0.0011135857
      10'd899: inv_x_count_prev = 16'b0000000001001001; // 1/899 = 0.0011123471
      10'd900: inv_x_count_prev = 16'b0000000001001001; // 1/900 = 0.0011111111
      10'd901: inv_x_count_prev = 16'b0000000001001001; // 1/901 = 0.0011098779
      10'd902: inv_x_count_prev = 16'b0000000001001001; // 1/902 = 0.0011086475
      10'd903: inv_x_count_prev = 16'b0000000001001001; // 1/903 = 0.0011074197
      10'd904: inv_x_count_prev = 16'b0000000001001000; // 1/904 = 0.0011061947
      10'd905: inv_x_count_prev = 16'b0000000001001000; // 1/905 = 0.0011049724
      10'd906: inv_x_count_prev = 16'b0000000001001000; // 1/906 = 0.0011037528
      10'd907: inv_x_count_prev = 16'b0000000001001000; // 1/907 = 0.0011025358
      10'd908: inv_x_count_prev = 16'b0000000001001000; // 1/908 = 0.0011013216
      10'd909: inv_x_count_prev = 16'b0000000001001000; // 1/909 = 0.0011001100
      10'd910: inv_x_count_prev = 16'b0000000001001000; // 1/910 = 0.0010989011
      10'd911: inv_x_count_prev = 16'b0000000001001000; // 1/911 = 0.0010976948
      10'd912: inv_x_count_prev = 16'b0000000001001000; // 1/912 = 0.0010964912
      10'd913: inv_x_count_prev = 16'b0000000001001000; // 1/913 = 0.0010952903
      10'd914: inv_x_count_prev = 16'b0000000001001000; // 1/914 = 0.0010940919
      10'd915: inv_x_count_prev = 16'b0000000001001000; // 1/915 = 0.0010928962
      10'd916: inv_x_count_prev = 16'b0000000001001000; // 1/916 = 0.0010917031
      10'd917: inv_x_count_prev = 16'b0000000001000111; // 1/917 = 0.0010905125
      10'd918: inv_x_count_prev = 16'b0000000001000111; // 1/918 = 0.0010893246
      10'd919: inv_x_count_prev = 16'b0000000001000111; // 1/919 = 0.0010881393
      10'd920: inv_x_count_prev = 16'b0000000001000111; // 1/920 = 0.0010869565
      10'd921: inv_x_count_prev = 16'b0000000001000111; // 1/921 = 0.0010857763
      10'd922: inv_x_count_prev = 16'b0000000001000111; // 1/922 = 0.0010845987
      10'd923: inv_x_count_prev = 16'b0000000001000111; // 1/923 = 0.0010834236
      10'd924: inv_x_count_prev = 16'b0000000001000111; // 1/924 = 0.0010822511
      10'd925: inv_x_count_prev = 16'b0000000001000111; // 1/925 = 0.0010810811
      10'd926: inv_x_count_prev = 16'b0000000001000111; // 1/926 = 0.0010799136
      10'd927: inv_x_count_prev = 16'b0000000001000111; // 1/927 = 0.0010787487
      10'd928: inv_x_count_prev = 16'b0000000001000111; // 1/928 = 0.0010775862
      10'd929: inv_x_count_prev = 16'b0000000001000111; // 1/929 = 0.0010764263
      10'd930: inv_x_count_prev = 16'b0000000001000110; // 1/930 = 0.0010752688
      10'd931: inv_x_count_prev = 16'b0000000001000110; // 1/931 = 0.0010741139
      10'd932: inv_x_count_prev = 16'b0000000001000110; // 1/932 = 0.0010729614
      10'd933: inv_x_count_prev = 16'b0000000001000110; // 1/933 = 0.0010718114
      10'd934: inv_x_count_prev = 16'b0000000001000110; // 1/934 = 0.0010706638
      10'd935: inv_x_count_prev = 16'b0000000001000110; // 1/935 = 0.0010695187
      10'd936: inv_x_count_prev = 16'b0000000001000110; // 1/936 = 0.0010683761
      10'd937: inv_x_count_prev = 16'b0000000001000110; // 1/937 = 0.0010672359
      10'd938: inv_x_count_prev = 16'b0000000001000110; // 1/938 = 0.0010660981
      10'd939: inv_x_count_prev = 16'b0000000001000110; // 1/939 = 0.0010649627
      10'd940: inv_x_count_prev = 16'b0000000001000110; // 1/940 = 0.0010638298
      10'd941: inv_x_count_prev = 16'b0000000001000110; // 1/941 = 0.0010626993
      10'd942: inv_x_count_prev = 16'b0000000001000110; // 1/942 = 0.0010615711
      10'd943: inv_x_count_prev = 16'b0000000001000101; // 1/943 = 0.0010604454
      10'd944: inv_x_count_prev = 16'b0000000001000101; // 1/944 = 0.0010593220
      10'd945: inv_x_count_prev = 16'b0000000001000101; // 1/945 = 0.0010582011
      10'd946: inv_x_count_prev = 16'b0000000001000101; // 1/946 = 0.0010570825
      10'd947: inv_x_count_prev = 16'b0000000001000101; // 1/947 = 0.0010559662
      10'd948: inv_x_count_prev = 16'b0000000001000101; // 1/948 = 0.0010548523
      10'd949: inv_x_count_prev = 16'b0000000001000101; // 1/949 = 0.0010537408
      10'd950: inv_x_count_prev = 16'b0000000001000101; // 1/950 = 0.0010526316
      10'd951: inv_x_count_prev = 16'b0000000001000101; // 1/951 = 0.0010515247
      10'd952: inv_x_count_prev = 16'b0000000001000101; // 1/952 = 0.0010504202
      10'd953: inv_x_count_prev = 16'b0000000001000101; // 1/953 = 0.0010493179
      10'd954: inv_x_count_prev = 16'b0000000001000101; // 1/954 = 0.0010482180
      10'd955: inv_x_count_prev = 16'b0000000001000101; // 1/955 = 0.0010471204
      10'd956: inv_x_count_prev = 16'b0000000001000101; // 1/956 = 0.0010460251
      10'd957: inv_x_count_prev = 16'b0000000001000100; // 1/957 = 0.0010449321
      10'd958: inv_x_count_prev = 16'b0000000001000100; // 1/958 = 0.0010438413
      10'd959: inv_x_count_prev = 16'b0000000001000100; // 1/959 = 0.0010427529
      10'd960: inv_x_count_prev = 16'b0000000001000100; // 1/960 = 0.0010416667
      10'd961: inv_x_count_prev = 16'b0000000001000100; // 1/961 = 0.0010405827
      10'd962: inv_x_count_prev = 16'b0000000001000100; // 1/962 = 0.0010395010
      10'd963: inv_x_count_prev = 16'b0000000001000100; // 1/963 = 0.0010384216
      10'd964: inv_x_count_prev = 16'b0000000001000100; // 1/964 = 0.0010373444
      10'd965: inv_x_count_prev = 16'b0000000001000100; // 1/965 = 0.0010362694
      10'd966: inv_x_count_prev = 16'b0000000001000100; // 1/966 = 0.0010351967
      10'd967: inv_x_count_prev = 16'b0000000001000100; // 1/967 = 0.0010341262
      10'd968: inv_x_count_prev = 16'b0000000001000100; // 1/968 = 0.0010330579
      10'd969: inv_x_count_prev = 16'b0000000001000100; // 1/969 = 0.0010319917
      10'd970: inv_x_count_prev = 16'b0000000001000100; // 1/970 = 0.0010309278
      10'd971: inv_x_count_prev = 16'b0000000001000011; // 1/971 = 0.0010298661
      10'd972: inv_x_count_prev = 16'b0000000001000011; // 1/972 = 0.0010288066
      10'd973: inv_x_count_prev = 16'b0000000001000011; // 1/973 = 0.0010277492
      10'd974: inv_x_count_prev = 16'b0000000001000011; // 1/974 = 0.0010266940
      10'd975: inv_x_count_prev = 16'b0000000001000011; // 1/975 = 0.0010256410
      10'd976: inv_x_count_prev = 16'b0000000001000011; // 1/976 = 0.0010245902
      10'd977: inv_x_count_prev = 16'b0000000001000011; // 1/977 = 0.0010235415
      10'd978: inv_x_count_prev = 16'b0000000001000011; // 1/978 = 0.0010224949
      10'd979: inv_x_count_prev = 16'b0000000001000011; // 1/979 = 0.0010214505
      10'd980: inv_x_count_prev = 16'b0000000001000011; // 1/980 = 0.0010204082
      10'd981: inv_x_count_prev = 16'b0000000001000011; // 1/981 = 0.0010193680
      10'd982: inv_x_count_prev = 16'b0000000001000011; // 1/982 = 0.0010183299
      10'd983: inv_x_count_prev = 16'b0000000001000011; // 1/983 = 0.0010172940
      10'd984: inv_x_count_prev = 16'b0000000001000011; // 1/984 = 0.0010162602
      10'd985: inv_x_count_prev = 16'b0000000001000011; // 1/985 = 0.0010152284
      10'd986: inv_x_count_prev = 16'b0000000001000010; // 1/986 = 0.0010141988
      10'd987: inv_x_count_prev = 16'b0000000001000010; // 1/987 = 0.0010131712
      10'd988: inv_x_count_prev = 16'b0000000001000010; // 1/988 = 0.0010121457
      10'd989: inv_x_count_prev = 16'b0000000001000010; // 1/989 = 0.0010111223
      10'd990: inv_x_count_prev = 16'b0000000001000010; // 1/990 = 0.0010101010
      10'd991: inv_x_count_prev = 16'b0000000001000010; // 1/991 = 0.0010090817
      10'd992: inv_x_count_prev = 16'b0000000001000010; // 1/992 = 0.0010080645
      10'd993: inv_x_count_prev = 16'b0000000001000010; // 1/993 = 0.0010070493
      10'd994: inv_x_count_prev = 16'b0000000001000010; // 1/994 = 0.0010060362
      10'd995: inv_x_count_prev = 16'b0000000001000010; // 1/995 = 0.0010050251
      10'd996: inv_x_count_prev = 16'b0000000001000010; // 1/996 = 0.0010040161
      10'd997: inv_x_count_prev = 16'b0000000001000010; // 1/997 = 0.0010030090
      10'd998: inv_x_count_prev = 16'b0000000001000010; // 1/998 = 0.0010020040
      10'd999: inv_x_count_prev = 16'b0000000001000010; // 1/999 = 0.0010010010
      10'd1000: inv_x_count_prev = 16'b0000000001000010; // 1/1000 = 0.0010000000
      10'd1001: inv_x_count_prev = 16'b0000000001000001; // 1/1001 = 0.0009990010
      10'd1002: inv_x_count_prev = 16'b0000000001000001; // 1/1002 = 0.0009980040
      10'd1003: inv_x_count_prev = 16'b0000000001000001; // 1/1003 = 0.0009970090
      10'd1004: inv_x_count_prev = 16'b0000000001000001; // 1/1004 = 0.0009960159
      10'd1005: inv_x_count_prev = 16'b0000000001000001; // 1/1005 = 0.0009950249
      10'd1006: inv_x_count_prev = 16'b0000000001000001; // 1/1006 = 0.0009940358
      10'd1007: inv_x_count_prev = 16'b0000000001000001; // 1/1007 = 0.0009930487
      10'd1008: inv_x_count_prev = 16'b0000000001000001; // 1/1008 = 0.0009920635
      10'd1009: inv_x_count_prev = 16'b0000000001000001; // 1/1009 = 0.0009910803
      10'd1010: inv_x_count_prev = 16'b0000000001000001; // 1/1010 = 0.0009900990
      10'd1011: inv_x_count_prev = 16'b0000000001000001; // 1/1011 = 0.0009891197
      10'd1012: inv_x_count_prev = 16'b0000000001000001; // 1/1012 = 0.0009881423
      10'd1013: inv_x_count_prev = 16'b0000000001000001; // 1/1013 = 0.0009871668
      10'd1014: inv_x_count_prev = 16'b0000000001000001; // 1/1014 = 0.0009861933
      10'd1015: inv_x_count_prev = 16'b0000000001000001; // 1/1015 = 0.0009852217
      10'd1016: inv_x_count_prev = 16'b0000000001000001; // 1/1016 = 0.0009842520
      10'd1017: inv_x_count_prev = 16'b0000000001000000; // 1/1017 = 0.0009832842
      10'd1018: inv_x_count_prev = 16'b0000000001000000; // 1/1018 = 0.0009823183
      10'd1019: inv_x_count_prev = 16'b0000000001000000; // 1/1019 = 0.0009813543
      10'd1020: inv_x_count_prev = 16'b0000000001000000; // 1/1020 = 0.0009803922
      10'd1021: inv_x_count_prev = 16'b0000000001000000; // 1/1021 = 0.0009794319
      10'd1022: inv_x_count_prev = 16'b0000000001000000; // 1/1022 = 0.0009784736
      10'd1023: inv_x_count_prev = 16'b0000000001000000; // 1/1023 = 0.0009775171
      10'd1024: inv_x_count_prev = 16'b0000000001000000; // 1/1024 = 0.0009765625
      default: inv_x_count_prev = '0; // Default case
    endcase
  end
//  always_comb begin
//    case (x_count+1)
//      10'd2: inv_x_count_next = 16'b1000000000000000; // 1/2 = 0.5000000000
//      10'd3: inv_x_count_next = 16'b0101010101010101; // 1/3 = 0.3333333333
//      10'd4: inv_x_count_next = 16'b0100000000000000; // 1/4 = 0.2500000000
//      10'd5: inv_x_count_next = 16'b0011001100110011; // 1/5 = 0.2000000000
//      10'd6: inv_x_count_next = 16'b0010101010101011; // 1/6 = 0.1666666667
//      10'd7: inv_x_count_next = 16'b0010010010010010; // 1/7 = 0.1428571429
//      10'd8: inv_x_count_next = 16'b0010000000000000; // 1/8 = 0.1250000000
//      10'd9: inv_x_count_next = 16'b0001110001110010; // 1/9 = 0.1111111111
//      10'd10: inv_x_count_next = 16'b0001100110011010; // 1/10 = 0.1000000000
//      10'd11: inv_x_count_next = 16'b0001011101000110; // 1/11 = 0.0909090909
//      10'd12: inv_x_count_next = 16'b0001010101010101; // 1/12 = 0.0833333333
//      10'd13: inv_x_count_next = 16'b0001001110110001; // 1/13 = 0.0769230769
//      10'd14: inv_x_count_next = 16'b0001001001001001; // 1/14 = 0.0714285714
//      10'd15: inv_x_count_next = 16'b0001000100010001; // 1/15 = 0.0666666667
//      10'd16: inv_x_count_next = 16'b0001000000000000; // 1/16 = 0.0625000000
//      10'd17: inv_x_count_next = 16'b0000111100001111; // 1/17 = 0.0588235294
//      10'd18: inv_x_count_next = 16'b0000111000111001; // 1/18 = 0.0555555556
//      10'd19: inv_x_count_next = 16'b0000110101111001; // 1/19 = 0.0526315789
//      10'd20: inv_x_count_next = 16'b0000110011001101; // 1/20 = 0.0500000000
//      10'd21: inv_x_count_next = 16'b0000110000110001; // 1/21 = 0.0476190476
//      10'd22: inv_x_count_next = 16'b0000101110100011; // 1/22 = 0.0454545455
//      10'd23: inv_x_count_next = 16'b0000101100100001; // 1/23 = 0.0434782609
//      10'd24: inv_x_count_next = 16'b0000101010101011; // 1/24 = 0.0416666667
//      10'd25: inv_x_count_next = 16'b0000101000111101; // 1/25 = 0.0400000000
//      10'd26: inv_x_count_next = 16'b0000100111011001; // 1/26 = 0.0384615385
//      10'd27: inv_x_count_next = 16'b0000100101111011; // 1/27 = 0.0370370370
//      10'd28: inv_x_count_next = 16'b0000100100100101; // 1/28 = 0.0357142857
//      10'd29: inv_x_count_next = 16'b0000100011010100; // 1/29 = 0.0344827586
//      10'd30: inv_x_count_next = 16'b0000100010001001; // 1/30 = 0.0333333333
//      10'd31: inv_x_count_next = 16'b0000100001000010; // 1/31 = 0.0322580645
//      10'd32: inv_x_count_next = 16'b0000100000000000; // 1/32 = 0.0312500000
//      10'd33: inv_x_count_next = 16'b0000011111000010; // 1/33 = 0.0303030303
//      10'd34: inv_x_count_next = 16'b0000011110001000; // 1/34 = 0.0294117647
//      10'd35: inv_x_count_next = 16'b0000011101010000; // 1/35 = 0.0285714286
//      10'd36: inv_x_count_next = 16'b0000011100011100; // 1/36 = 0.0277777778
//      10'd37: inv_x_count_next = 16'b0000011011101011; // 1/37 = 0.0270270270
//      10'd38: inv_x_count_next = 16'b0000011010111101; // 1/38 = 0.0263157895
//      10'd39: inv_x_count_next = 16'b0000011010010000; // 1/39 = 0.0256410256
//      10'd40: inv_x_count_next = 16'b0000011001100110; // 1/40 = 0.0250000000
//      10'd41: inv_x_count_next = 16'b0000011000111110; // 1/41 = 0.0243902439
//      10'd42: inv_x_count_next = 16'b0000011000011000; // 1/42 = 0.0238095238
//      10'd43: inv_x_count_next = 16'b0000010111110100; // 1/43 = 0.0232558140
//      10'd44: inv_x_count_next = 16'b0000010111010001; // 1/44 = 0.0227272727
//      10'd45: inv_x_count_next = 16'b0000010110110000; // 1/45 = 0.0222222222
//      10'd46: inv_x_count_next = 16'b0000010110010001; // 1/46 = 0.0217391304
//      10'd47: inv_x_count_next = 16'b0000010101110010; // 1/47 = 0.0212765957
//      10'd48: inv_x_count_next = 16'b0000010101010101; // 1/48 = 0.0208333333
//      10'd49: inv_x_count_next = 16'b0000010100111001; // 1/49 = 0.0204081633
//      10'd50: inv_x_count_next = 16'b0000010100011111; // 1/50 = 0.0200000000
//      10'd51: inv_x_count_next = 16'b0000010100000101; // 1/51 = 0.0196078431
//      10'd52: inv_x_count_next = 16'b0000010011101100; // 1/52 = 0.0192307692
//      10'd53: inv_x_count_next = 16'b0000010011010101; // 1/53 = 0.0188679245
//      10'd54: inv_x_count_next = 16'b0000010010111110; // 1/54 = 0.0185185185
//      10'd55: inv_x_count_next = 16'b0000010010101000; // 1/55 = 0.0181818182
//      10'd56: inv_x_count_next = 16'b0000010010010010; // 1/56 = 0.0178571429
//      10'd57: inv_x_count_next = 16'b0000010001111110; // 1/57 = 0.0175438596
//      10'd58: inv_x_count_next = 16'b0000010001101010; // 1/58 = 0.0172413793
//      10'd59: inv_x_count_next = 16'b0000010001010111; // 1/59 = 0.0169491525
//      10'd60: inv_x_count_next = 16'b0000010001000100; // 1/60 = 0.0166666667
//      10'd61: inv_x_count_next = 16'b0000010000110010; // 1/61 = 0.0163934426
//      10'd62: inv_x_count_next = 16'b0000010000100001; // 1/62 = 0.0161290323
//      10'd63: inv_x_count_next = 16'b0000010000010000; // 1/63 = 0.0158730159
//      10'd64: inv_x_count_next = 16'b0000010000000000; // 1/64 = 0.0156250000
//      10'd65: inv_x_count_next = 16'b0000001111110000; // 1/65 = 0.0153846154
//      10'd66: inv_x_count_next = 16'b0000001111100001; // 1/66 = 0.0151515152
//      10'd67: inv_x_count_next = 16'b0000001111010010; // 1/67 = 0.0149253731
//      10'd68: inv_x_count_next = 16'b0000001111000100; // 1/68 = 0.0147058824
//      10'd69: inv_x_count_next = 16'b0000001110110110; // 1/69 = 0.0144927536
//      10'd70: inv_x_count_next = 16'b0000001110101000; // 1/70 = 0.0142857143
//      10'd71: inv_x_count_next = 16'b0000001110011011; // 1/71 = 0.0140845070
//      10'd72: inv_x_count_next = 16'b0000001110001110; // 1/72 = 0.0138888889
//      10'd73: inv_x_count_next = 16'b0000001110000010; // 1/73 = 0.0136986301
//      10'd74: inv_x_count_next = 16'b0000001101110110; // 1/74 = 0.0135135135
//      10'd75: inv_x_count_next = 16'b0000001101101010; // 1/75 = 0.0133333333
//      10'd76: inv_x_count_next = 16'b0000001101011110; // 1/76 = 0.0131578947
//      10'd77: inv_x_count_next = 16'b0000001101010011; // 1/77 = 0.0129870130
//      10'd78: inv_x_count_next = 16'b0000001101001000; // 1/78 = 0.0128205128
//      10'd79: inv_x_count_next = 16'b0000001100111110; // 1/79 = 0.0126582278
//      10'd80: inv_x_count_next = 16'b0000001100110011; // 1/80 = 0.0125000000
//      10'd81: inv_x_count_next = 16'b0000001100101001; // 1/81 = 0.0123456790
//      10'd82: inv_x_count_next = 16'b0000001100011111; // 1/82 = 0.0121951220
//      10'd83: inv_x_count_next = 16'b0000001100010110; // 1/83 = 0.0120481928
//      10'd84: inv_x_count_next = 16'b0000001100001100; // 1/84 = 0.0119047619
//      10'd85: inv_x_count_next = 16'b0000001100000011; // 1/85 = 0.0117647059
//      10'd86: inv_x_count_next = 16'b0000001011111010; // 1/86 = 0.0116279070
//      10'd87: inv_x_count_next = 16'b0000001011110001; // 1/87 = 0.0114942529
//      10'd88: inv_x_count_next = 16'b0000001011101001; // 1/88 = 0.0113636364
//      10'd89: inv_x_count_next = 16'b0000001011100000; // 1/89 = 0.0112359551
//      10'd90: inv_x_count_next = 16'b0000001011011000; // 1/90 = 0.0111111111
//      10'd91: inv_x_count_next = 16'b0000001011010000; // 1/91 = 0.0109890110
//      10'd92: inv_x_count_next = 16'b0000001011001000; // 1/92 = 0.0108695652
//      10'd93: inv_x_count_next = 16'b0000001011000001; // 1/93 = 0.0107526882
//      10'd94: inv_x_count_next = 16'b0000001010111001; // 1/94 = 0.0106382979
//      10'd95: inv_x_count_next = 16'b0000001010110010; // 1/95 = 0.0105263158
//      10'd96: inv_x_count_next = 16'b0000001010101011; // 1/96 = 0.0104166667
//      10'd97: inv_x_count_next = 16'b0000001010100100; // 1/97 = 0.0103092784
//      10'd98: inv_x_count_next = 16'b0000001010011101; // 1/98 = 0.0102040816
//      10'd99: inv_x_count_next = 16'b0000001010010110; // 1/99 = 0.0101010101
//      10'd100: inv_x_count_next = 16'b0000001010001111; // 1/100 = 0.0100000000
//      10'd101: inv_x_count_next = 16'b0000001010001001; // 1/101 = 0.0099009901
//      10'd102: inv_x_count_next = 16'b0000001010000011; // 1/102 = 0.0098039216
//      10'd103: inv_x_count_next = 16'b0000001001111100; // 1/103 = 0.0097087379
//      10'd104: inv_x_count_next = 16'b0000001001110110; // 1/104 = 0.0096153846
//      10'd105: inv_x_count_next = 16'b0000001001110000; // 1/105 = 0.0095238095
//      10'd106: inv_x_count_next = 16'b0000001001101010; // 1/106 = 0.0094339623
//      10'd107: inv_x_count_next = 16'b0000001001100100; // 1/107 = 0.0093457944
//      10'd108: inv_x_count_next = 16'b0000001001011111; // 1/108 = 0.0092592593
//      10'd109: inv_x_count_next = 16'b0000001001011001; // 1/109 = 0.0091743119
//      10'd110: inv_x_count_next = 16'b0000001001010100; // 1/110 = 0.0090909091
//      10'd111: inv_x_count_next = 16'b0000001001001110; // 1/111 = 0.0090090090
//      10'd112: inv_x_count_next = 16'b0000001001001001; // 1/112 = 0.0089285714
//      10'd113: inv_x_count_next = 16'b0000001001000100; // 1/113 = 0.0088495575
//      10'd114: inv_x_count_next = 16'b0000001000111111; // 1/114 = 0.0087719298
//      10'd115: inv_x_count_next = 16'b0000001000111010; // 1/115 = 0.0086956522
//      10'd116: inv_x_count_next = 16'b0000001000110101; // 1/116 = 0.0086206897
//      10'd117: inv_x_count_next = 16'b0000001000110000; // 1/117 = 0.0085470085
//      10'd118: inv_x_count_next = 16'b0000001000101011; // 1/118 = 0.0084745763
//      10'd119: inv_x_count_next = 16'b0000001000100111; // 1/119 = 0.0084033613
//      10'd120: inv_x_count_next = 16'b0000001000100010; // 1/120 = 0.0083333333
//      10'd121: inv_x_count_next = 16'b0000001000011110; // 1/121 = 0.0082644628
//      10'd122: inv_x_count_next = 16'b0000001000011001; // 1/122 = 0.0081967213
//      10'd123: inv_x_count_next = 16'b0000001000010101; // 1/123 = 0.0081300813
//      10'd124: inv_x_count_next = 16'b0000001000010001; // 1/124 = 0.0080645161
//      10'd125: inv_x_count_next = 16'b0000001000001100; // 1/125 = 0.0080000000
//      10'd126: inv_x_count_next = 16'b0000001000001000; // 1/126 = 0.0079365079
//      10'd127: inv_x_count_next = 16'b0000001000000100; // 1/127 = 0.0078740157
//      10'd128: inv_x_count_next = 16'b0000001000000000; // 1/128 = 0.0078125000
//      10'd129: inv_x_count_next = 16'b0000000111111100; // 1/129 = 0.0077519380
//      10'd130: inv_x_count_next = 16'b0000000111111000; // 1/130 = 0.0076923077
//      10'd131: inv_x_count_next = 16'b0000000111110100; // 1/131 = 0.0076335878
//      10'd132: inv_x_count_next = 16'b0000000111110000; // 1/132 = 0.0075757576
//      10'd133: inv_x_count_next = 16'b0000000111101101; // 1/133 = 0.0075187970
//      10'd134: inv_x_count_next = 16'b0000000111101001; // 1/134 = 0.0074626866
//      10'd135: inv_x_count_next = 16'b0000000111100101; // 1/135 = 0.0074074074
//      10'd136: inv_x_count_next = 16'b0000000111100010; // 1/136 = 0.0073529412
//      10'd137: inv_x_count_next = 16'b0000000111011110; // 1/137 = 0.0072992701
//      10'd138: inv_x_count_next = 16'b0000000111011011; // 1/138 = 0.0072463768
//      10'd139: inv_x_count_next = 16'b0000000111010111; // 1/139 = 0.0071942446
//      10'd140: inv_x_count_next = 16'b0000000111010100; // 1/140 = 0.0071428571
//      10'd141: inv_x_count_next = 16'b0000000111010001; // 1/141 = 0.0070921986
//      10'd142: inv_x_count_next = 16'b0000000111001110; // 1/142 = 0.0070422535
//      10'd143: inv_x_count_next = 16'b0000000111001010; // 1/143 = 0.0069930070
//      10'd144: inv_x_count_next = 16'b0000000111000111; // 1/144 = 0.0069444444
//      10'd145: inv_x_count_next = 16'b0000000111000100; // 1/145 = 0.0068965517
//      10'd146: inv_x_count_next = 16'b0000000111000001; // 1/146 = 0.0068493151
//      10'd147: inv_x_count_next = 16'b0000000110111110; // 1/147 = 0.0068027211
//      10'd148: inv_x_count_next = 16'b0000000110111011; // 1/148 = 0.0067567568
//      10'd149: inv_x_count_next = 16'b0000000110111000; // 1/149 = 0.0067114094
//      10'd150: inv_x_count_next = 16'b0000000110110101; // 1/150 = 0.0066666667
//      10'd151: inv_x_count_next = 16'b0000000110110010; // 1/151 = 0.0066225166
//      10'd152: inv_x_count_next = 16'b0000000110101111; // 1/152 = 0.0065789474
//      10'd153: inv_x_count_next = 16'b0000000110101100; // 1/153 = 0.0065359477
//      10'd154: inv_x_count_next = 16'b0000000110101010; // 1/154 = 0.0064935065
//      10'd155: inv_x_count_next = 16'b0000000110100111; // 1/155 = 0.0064516129
//      10'd156: inv_x_count_next = 16'b0000000110100100; // 1/156 = 0.0064102564
//      10'd157: inv_x_count_next = 16'b0000000110100001; // 1/157 = 0.0063694268
//      10'd158: inv_x_count_next = 16'b0000000110011111; // 1/158 = 0.0063291139
//      10'd159: inv_x_count_next = 16'b0000000110011100; // 1/159 = 0.0062893082
//      10'd160: inv_x_count_next = 16'b0000000110011010; // 1/160 = 0.0062500000
//      10'd161: inv_x_count_next = 16'b0000000110010111; // 1/161 = 0.0062111801
//      10'd162: inv_x_count_next = 16'b0000000110010101; // 1/162 = 0.0061728395
//      10'd163: inv_x_count_next = 16'b0000000110010010; // 1/163 = 0.0061349693
//      10'd164: inv_x_count_next = 16'b0000000110010000; // 1/164 = 0.0060975610
//      10'd165: inv_x_count_next = 16'b0000000110001101; // 1/165 = 0.0060606061
//      10'd166: inv_x_count_next = 16'b0000000110001011; // 1/166 = 0.0060240964
//      10'd167: inv_x_count_next = 16'b0000000110001000; // 1/167 = 0.0059880240
//      10'd168: inv_x_count_next = 16'b0000000110000110; // 1/168 = 0.0059523810
//      10'd169: inv_x_count_next = 16'b0000000110000100; // 1/169 = 0.0059171598
//      10'd170: inv_x_count_next = 16'b0000000110000010; // 1/170 = 0.0058823529
//      10'd171: inv_x_count_next = 16'b0000000101111111; // 1/171 = 0.0058479532
//      10'd172: inv_x_count_next = 16'b0000000101111101; // 1/172 = 0.0058139535
//      10'd173: inv_x_count_next = 16'b0000000101111011; // 1/173 = 0.0057803468
//      10'd174: inv_x_count_next = 16'b0000000101111001; // 1/174 = 0.0057471264
//      10'd175: inv_x_count_next = 16'b0000000101110110; // 1/175 = 0.0057142857
//      10'd176: inv_x_count_next = 16'b0000000101110100; // 1/176 = 0.0056818182
//      10'd177: inv_x_count_next = 16'b0000000101110010; // 1/177 = 0.0056497175
//      10'd178: inv_x_count_next = 16'b0000000101110000; // 1/178 = 0.0056179775
//      10'd179: inv_x_count_next = 16'b0000000101101110; // 1/179 = 0.0055865922
//      10'd180: inv_x_count_next = 16'b0000000101101100; // 1/180 = 0.0055555556
//      10'd181: inv_x_count_next = 16'b0000000101101010; // 1/181 = 0.0055248619
//      10'd182: inv_x_count_next = 16'b0000000101101000; // 1/182 = 0.0054945055
//      10'd183: inv_x_count_next = 16'b0000000101100110; // 1/183 = 0.0054644809
//      10'd184: inv_x_count_next = 16'b0000000101100100; // 1/184 = 0.0054347826
//      10'd185: inv_x_count_next = 16'b0000000101100010; // 1/185 = 0.0054054054
//      10'd186: inv_x_count_next = 16'b0000000101100000; // 1/186 = 0.0053763441
//      10'd187: inv_x_count_next = 16'b0000000101011110; // 1/187 = 0.0053475936
//      10'd188: inv_x_count_next = 16'b0000000101011101; // 1/188 = 0.0053191489
//      10'd189: inv_x_count_next = 16'b0000000101011011; // 1/189 = 0.0052910053
//      10'd190: inv_x_count_next = 16'b0000000101011001; // 1/190 = 0.0052631579
//      10'd191: inv_x_count_next = 16'b0000000101010111; // 1/191 = 0.0052356021
//      10'd192: inv_x_count_next = 16'b0000000101010101; // 1/192 = 0.0052083333
//      10'd193: inv_x_count_next = 16'b0000000101010100; // 1/193 = 0.0051813472
//      10'd194: inv_x_count_next = 16'b0000000101010010; // 1/194 = 0.0051546392
//      10'd195: inv_x_count_next = 16'b0000000101010000; // 1/195 = 0.0051282051
//      10'd196: inv_x_count_next = 16'b0000000101001110; // 1/196 = 0.0051020408
//      10'd197: inv_x_count_next = 16'b0000000101001101; // 1/197 = 0.0050761421
//      10'd198: inv_x_count_next = 16'b0000000101001011; // 1/198 = 0.0050505051
//      10'd199: inv_x_count_next = 16'b0000000101001001; // 1/199 = 0.0050251256
//      10'd200: inv_x_count_next = 16'b0000000101001000; // 1/200 = 0.0050000000
//      10'd201: inv_x_count_next = 16'b0000000101000110; // 1/201 = 0.0049751244
//      10'd202: inv_x_count_next = 16'b0000000101000100; // 1/202 = 0.0049504950
//      10'd203: inv_x_count_next = 16'b0000000101000011; // 1/203 = 0.0049261084
//      10'd204: inv_x_count_next = 16'b0000000101000001; // 1/204 = 0.0049019608
//      10'd205: inv_x_count_next = 16'b0000000101000000; // 1/205 = 0.0048780488
//      10'd206: inv_x_count_next = 16'b0000000100111110; // 1/206 = 0.0048543689
//      10'd207: inv_x_count_next = 16'b0000000100111101; // 1/207 = 0.0048309179
//      10'd208: inv_x_count_next = 16'b0000000100111011; // 1/208 = 0.0048076923
//      10'd209: inv_x_count_next = 16'b0000000100111010; // 1/209 = 0.0047846890
//      10'd210: inv_x_count_next = 16'b0000000100111000; // 1/210 = 0.0047619048
//      10'd211: inv_x_count_next = 16'b0000000100110111; // 1/211 = 0.0047393365
//      10'd212: inv_x_count_next = 16'b0000000100110101; // 1/212 = 0.0047169811
//      10'd213: inv_x_count_next = 16'b0000000100110100; // 1/213 = 0.0046948357
//      10'd214: inv_x_count_next = 16'b0000000100110010; // 1/214 = 0.0046728972
//      10'd215: inv_x_count_next = 16'b0000000100110001; // 1/215 = 0.0046511628
//      10'd216: inv_x_count_next = 16'b0000000100101111; // 1/216 = 0.0046296296
//      10'd217: inv_x_count_next = 16'b0000000100101110; // 1/217 = 0.0046082949
//      10'd218: inv_x_count_next = 16'b0000000100101101; // 1/218 = 0.0045871560
//      10'd219: inv_x_count_next = 16'b0000000100101011; // 1/219 = 0.0045662100
//      10'd220: inv_x_count_next = 16'b0000000100101010; // 1/220 = 0.0045454545
//      10'd221: inv_x_count_next = 16'b0000000100101001; // 1/221 = 0.0045248869
//      10'd222: inv_x_count_next = 16'b0000000100100111; // 1/222 = 0.0045045045
//      10'd223: inv_x_count_next = 16'b0000000100100110; // 1/223 = 0.0044843049
//      10'd224: inv_x_count_next = 16'b0000000100100101; // 1/224 = 0.0044642857
//      10'd225: inv_x_count_next = 16'b0000000100100011; // 1/225 = 0.0044444444
//      10'd226: inv_x_count_next = 16'b0000000100100010; // 1/226 = 0.0044247788
//      10'd227: inv_x_count_next = 16'b0000000100100001; // 1/227 = 0.0044052863
//      10'd228: inv_x_count_next = 16'b0000000100011111; // 1/228 = 0.0043859649
//      10'd229: inv_x_count_next = 16'b0000000100011110; // 1/229 = 0.0043668122
//      10'd230: inv_x_count_next = 16'b0000000100011101; // 1/230 = 0.0043478261
//      10'd231: inv_x_count_next = 16'b0000000100011100; // 1/231 = 0.0043290043
//      10'd232: inv_x_count_next = 16'b0000000100011010; // 1/232 = 0.0043103448
//      10'd233: inv_x_count_next = 16'b0000000100011001; // 1/233 = 0.0042918455
//      10'd234: inv_x_count_next = 16'b0000000100011000; // 1/234 = 0.0042735043
//      10'd235: inv_x_count_next = 16'b0000000100010111; // 1/235 = 0.0042553191
//      10'd236: inv_x_count_next = 16'b0000000100010110; // 1/236 = 0.0042372881
//      10'd237: inv_x_count_next = 16'b0000000100010101; // 1/237 = 0.0042194093
//      10'd238: inv_x_count_next = 16'b0000000100010011; // 1/238 = 0.0042016807
//      10'd239: inv_x_count_next = 16'b0000000100010010; // 1/239 = 0.0041841004
//      10'd240: inv_x_count_next = 16'b0000000100010001; // 1/240 = 0.0041666667
//      10'd241: inv_x_count_next = 16'b0000000100010000; // 1/241 = 0.0041493776
//      10'd242: inv_x_count_next = 16'b0000000100001111; // 1/242 = 0.0041322314
//      10'd243: inv_x_count_next = 16'b0000000100001110; // 1/243 = 0.0041152263
//      10'd244: inv_x_count_next = 16'b0000000100001101; // 1/244 = 0.0040983607
//      10'd245: inv_x_count_next = 16'b0000000100001011; // 1/245 = 0.0040816327
//      10'd246: inv_x_count_next = 16'b0000000100001010; // 1/246 = 0.0040650407
//      10'd247: inv_x_count_next = 16'b0000000100001001; // 1/247 = 0.0040485830
//      10'd248: inv_x_count_next = 16'b0000000100001000; // 1/248 = 0.0040322581
//      10'd249: inv_x_count_next = 16'b0000000100000111; // 1/249 = 0.0040160643
//      10'd250: inv_x_count_next = 16'b0000000100000110; // 1/250 = 0.0040000000
//      10'd251: inv_x_count_next = 16'b0000000100000101; // 1/251 = 0.0039840637
//      10'd252: inv_x_count_next = 16'b0000000100000100; // 1/252 = 0.0039682540
//      10'd253: inv_x_count_next = 16'b0000000100000011; // 1/253 = 0.0039525692
//      10'd254: inv_x_count_next = 16'b0000000100000010; // 1/254 = 0.0039370079
//      10'd255: inv_x_count_next = 16'b0000000100000001; // 1/255 = 0.0039215686
//      10'd256: inv_x_count_next = 16'b0000000100000000; // 1/256 = 0.0039062500
//      10'd257: inv_x_count_next = 16'b0000000011111111; // 1/257 = 0.0038910506
//      10'd258: inv_x_count_next = 16'b0000000011111110; // 1/258 = 0.0038759690
//      10'd259: inv_x_count_next = 16'b0000000011111101; // 1/259 = 0.0038610039
//      10'd260: inv_x_count_next = 16'b0000000011111100; // 1/260 = 0.0038461538
//      10'd261: inv_x_count_next = 16'b0000000011111011; // 1/261 = 0.0038314176
//      10'd262: inv_x_count_next = 16'b0000000011111010; // 1/262 = 0.0038167939
//      10'd263: inv_x_count_next = 16'b0000000011111001; // 1/263 = 0.0038022814
//      10'd264: inv_x_count_next = 16'b0000000011111000; // 1/264 = 0.0037878788
//      10'd265: inv_x_count_next = 16'b0000000011110111; // 1/265 = 0.0037735849
//      10'd266: inv_x_count_next = 16'b0000000011110110; // 1/266 = 0.0037593985
//      10'd267: inv_x_count_next = 16'b0000000011110101; // 1/267 = 0.0037453184
//      10'd268: inv_x_count_next = 16'b0000000011110101; // 1/268 = 0.0037313433
//      10'd269: inv_x_count_next = 16'b0000000011110100; // 1/269 = 0.0037174721
//      10'd270: inv_x_count_next = 16'b0000000011110011; // 1/270 = 0.0037037037
//      10'd271: inv_x_count_next = 16'b0000000011110010; // 1/271 = 0.0036900369
//      10'd272: inv_x_count_next = 16'b0000000011110001; // 1/272 = 0.0036764706
//      10'd273: inv_x_count_next = 16'b0000000011110000; // 1/273 = 0.0036630037
//      10'd274: inv_x_count_next = 16'b0000000011101111; // 1/274 = 0.0036496350
//      10'd275: inv_x_count_next = 16'b0000000011101110; // 1/275 = 0.0036363636
//      10'd276: inv_x_count_next = 16'b0000000011101101; // 1/276 = 0.0036231884
//      10'd277: inv_x_count_next = 16'b0000000011101101; // 1/277 = 0.0036101083
//      10'd278: inv_x_count_next = 16'b0000000011101100; // 1/278 = 0.0035971223
//      10'd279: inv_x_count_next = 16'b0000000011101011; // 1/279 = 0.0035842294
//      10'd280: inv_x_count_next = 16'b0000000011101010; // 1/280 = 0.0035714286
//      10'd281: inv_x_count_next = 16'b0000000011101001; // 1/281 = 0.0035587189
//      10'd282: inv_x_count_next = 16'b0000000011101000; // 1/282 = 0.0035460993
//      10'd283: inv_x_count_next = 16'b0000000011101000; // 1/283 = 0.0035335689
//      10'd284: inv_x_count_next = 16'b0000000011100111; // 1/284 = 0.0035211268
//      10'd285: inv_x_count_next = 16'b0000000011100110; // 1/285 = 0.0035087719
//      10'd286: inv_x_count_next = 16'b0000000011100101; // 1/286 = 0.0034965035
//      10'd287: inv_x_count_next = 16'b0000000011100100; // 1/287 = 0.0034843206
//      10'd288: inv_x_count_next = 16'b0000000011100100; // 1/288 = 0.0034722222
//      10'd289: inv_x_count_next = 16'b0000000011100011; // 1/289 = 0.0034602076
//      10'd290: inv_x_count_next = 16'b0000000011100010; // 1/290 = 0.0034482759
//      10'd291: inv_x_count_next = 16'b0000000011100001; // 1/291 = 0.0034364261
//      10'd292: inv_x_count_next = 16'b0000000011100000; // 1/292 = 0.0034246575
//      10'd293: inv_x_count_next = 16'b0000000011100000; // 1/293 = 0.0034129693
//      10'd294: inv_x_count_next = 16'b0000000011011111; // 1/294 = 0.0034013605
//      10'd295: inv_x_count_next = 16'b0000000011011110; // 1/295 = 0.0033898305
//      10'd296: inv_x_count_next = 16'b0000000011011101; // 1/296 = 0.0033783784
//      10'd297: inv_x_count_next = 16'b0000000011011101; // 1/297 = 0.0033670034
//      10'd298: inv_x_count_next = 16'b0000000011011100; // 1/298 = 0.0033557047
//      10'd299: inv_x_count_next = 16'b0000000011011011; // 1/299 = 0.0033444816
//      10'd300: inv_x_count_next = 16'b0000000011011010; // 1/300 = 0.0033333333
//      10'd301: inv_x_count_next = 16'b0000000011011010; // 1/301 = 0.0033222591
//      10'd302: inv_x_count_next = 16'b0000000011011001; // 1/302 = 0.0033112583
//      10'd303: inv_x_count_next = 16'b0000000011011000; // 1/303 = 0.0033003300
//      10'd304: inv_x_count_next = 16'b0000000011011000; // 1/304 = 0.0032894737
//      10'd305: inv_x_count_next = 16'b0000000011010111; // 1/305 = 0.0032786885
//      10'd306: inv_x_count_next = 16'b0000000011010110; // 1/306 = 0.0032679739
//      10'd307: inv_x_count_next = 16'b0000000011010101; // 1/307 = 0.0032573290
//      10'd308: inv_x_count_next = 16'b0000000011010101; // 1/308 = 0.0032467532
//      10'd309: inv_x_count_next = 16'b0000000011010100; // 1/309 = 0.0032362460
//      10'd310: inv_x_count_next = 16'b0000000011010011; // 1/310 = 0.0032258065
//      10'd311: inv_x_count_next = 16'b0000000011010011; // 1/311 = 0.0032154341
//      10'd312: inv_x_count_next = 16'b0000000011010010; // 1/312 = 0.0032051282
//      10'd313: inv_x_count_next = 16'b0000000011010001; // 1/313 = 0.0031948882
//      10'd314: inv_x_count_next = 16'b0000000011010001; // 1/314 = 0.0031847134
//      10'd315: inv_x_count_next = 16'b0000000011010000; // 1/315 = 0.0031746032
//      10'd316: inv_x_count_next = 16'b0000000011001111; // 1/316 = 0.0031645570
//      10'd317: inv_x_count_next = 16'b0000000011001111; // 1/317 = 0.0031545741
//      10'd318: inv_x_count_next = 16'b0000000011001110; // 1/318 = 0.0031446541
//      10'd319: inv_x_count_next = 16'b0000000011001101; // 1/319 = 0.0031347962
//      10'd320: inv_x_count_next = 16'b0000000011001101; // 1/320 = 0.0031250000
//      10'd321: inv_x_count_next = 16'b0000000011001100; // 1/321 = 0.0031152648
//      10'd322: inv_x_count_next = 16'b0000000011001100; // 1/322 = 0.0031055901
//      10'd323: inv_x_count_next = 16'b0000000011001011; // 1/323 = 0.0030959752
//      10'd324: inv_x_count_next = 16'b0000000011001010; // 1/324 = 0.0030864198
//      10'd325: inv_x_count_next = 16'b0000000011001010; // 1/325 = 0.0030769231
//      10'd326: inv_x_count_next = 16'b0000000011001001; // 1/326 = 0.0030674847
//      10'd327: inv_x_count_next = 16'b0000000011001000; // 1/327 = 0.0030581040
//      10'd328: inv_x_count_next = 16'b0000000011001000; // 1/328 = 0.0030487805
//      10'd329: inv_x_count_next = 16'b0000000011000111; // 1/329 = 0.0030395137
//      10'd330: inv_x_count_next = 16'b0000000011000111; // 1/330 = 0.0030303030
//      10'd331: inv_x_count_next = 16'b0000000011000110; // 1/331 = 0.0030211480
//      10'd332: inv_x_count_next = 16'b0000000011000101; // 1/332 = 0.0030120482
//      10'd333: inv_x_count_next = 16'b0000000011000101; // 1/333 = 0.0030030030
//      10'd334: inv_x_count_next = 16'b0000000011000100; // 1/334 = 0.0029940120
//      10'd335: inv_x_count_next = 16'b0000000011000100; // 1/335 = 0.0029850746
//      10'd336: inv_x_count_next = 16'b0000000011000011; // 1/336 = 0.0029761905
//      10'd337: inv_x_count_next = 16'b0000000011000010; // 1/337 = 0.0029673591
//      10'd338: inv_x_count_next = 16'b0000000011000010; // 1/338 = 0.0029585799
//      10'd339: inv_x_count_next = 16'b0000000011000001; // 1/339 = 0.0029498525
//      10'd340: inv_x_count_next = 16'b0000000011000001; // 1/340 = 0.0029411765
//      10'd341: inv_x_count_next = 16'b0000000011000000; // 1/341 = 0.0029325513
//      10'd342: inv_x_count_next = 16'b0000000011000000; // 1/342 = 0.0029239766
//      10'd343: inv_x_count_next = 16'b0000000010111111; // 1/343 = 0.0029154519
//      10'd344: inv_x_count_next = 16'b0000000010111111; // 1/344 = 0.0029069767
//      10'd345: inv_x_count_next = 16'b0000000010111110; // 1/345 = 0.0028985507
//      10'd346: inv_x_count_next = 16'b0000000010111101; // 1/346 = 0.0028901734
//      10'd347: inv_x_count_next = 16'b0000000010111101; // 1/347 = 0.0028818444
//      10'd348: inv_x_count_next = 16'b0000000010111100; // 1/348 = 0.0028735632
//      10'd349: inv_x_count_next = 16'b0000000010111100; // 1/349 = 0.0028653295
//      10'd350: inv_x_count_next = 16'b0000000010111011; // 1/350 = 0.0028571429
//      10'd351: inv_x_count_next = 16'b0000000010111011; // 1/351 = 0.0028490028
//      10'd352: inv_x_count_next = 16'b0000000010111010; // 1/352 = 0.0028409091
//      10'd353: inv_x_count_next = 16'b0000000010111010; // 1/353 = 0.0028328612
//      10'd354: inv_x_count_next = 16'b0000000010111001; // 1/354 = 0.0028248588
//      10'd355: inv_x_count_next = 16'b0000000010111001; // 1/355 = 0.0028169014
//      10'd356: inv_x_count_next = 16'b0000000010111000; // 1/356 = 0.0028089888
//      10'd357: inv_x_count_next = 16'b0000000010111000; // 1/357 = 0.0028011204
//      10'd358: inv_x_count_next = 16'b0000000010110111; // 1/358 = 0.0027932961
//      10'd359: inv_x_count_next = 16'b0000000010110111; // 1/359 = 0.0027855153
//      10'd360: inv_x_count_next = 16'b0000000010110110; // 1/360 = 0.0027777778
//      10'd361: inv_x_count_next = 16'b0000000010110110; // 1/361 = 0.0027700831
//      10'd362: inv_x_count_next = 16'b0000000010110101; // 1/362 = 0.0027624309
//      10'd363: inv_x_count_next = 16'b0000000010110101; // 1/363 = 0.0027548209
//      10'd364: inv_x_count_next = 16'b0000000010110100; // 1/364 = 0.0027472527
//      10'd365: inv_x_count_next = 16'b0000000010110100; // 1/365 = 0.0027397260
//      10'd366: inv_x_count_next = 16'b0000000010110011; // 1/366 = 0.0027322404
//      10'd367: inv_x_count_next = 16'b0000000010110011; // 1/367 = 0.0027247956
//      10'd368: inv_x_count_next = 16'b0000000010110010; // 1/368 = 0.0027173913
//      10'd369: inv_x_count_next = 16'b0000000010110010; // 1/369 = 0.0027100271
//      10'd370: inv_x_count_next = 16'b0000000010110001; // 1/370 = 0.0027027027
//      10'd371: inv_x_count_next = 16'b0000000010110001; // 1/371 = 0.0026954178
//      10'd372: inv_x_count_next = 16'b0000000010110000; // 1/372 = 0.0026881720
//      10'd373: inv_x_count_next = 16'b0000000010110000; // 1/373 = 0.0026809651
//      10'd374: inv_x_count_next = 16'b0000000010101111; // 1/374 = 0.0026737968
//      10'd375: inv_x_count_next = 16'b0000000010101111; // 1/375 = 0.0026666667
//      10'd376: inv_x_count_next = 16'b0000000010101110; // 1/376 = 0.0026595745
//      10'd377: inv_x_count_next = 16'b0000000010101110; // 1/377 = 0.0026525199
//      10'd378: inv_x_count_next = 16'b0000000010101101; // 1/378 = 0.0026455026
//      10'd379: inv_x_count_next = 16'b0000000010101101; // 1/379 = 0.0026385224
//      10'd380: inv_x_count_next = 16'b0000000010101100; // 1/380 = 0.0026315789
//      10'd381: inv_x_count_next = 16'b0000000010101100; // 1/381 = 0.0026246719
//      10'd382: inv_x_count_next = 16'b0000000010101100; // 1/382 = 0.0026178010
//      10'd383: inv_x_count_next = 16'b0000000010101011; // 1/383 = 0.0026109661
//      10'd384: inv_x_count_next = 16'b0000000010101011; // 1/384 = 0.0026041667
//      10'd385: inv_x_count_next = 16'b0000000010101010; // 1/385 = 0.0025974026
//      10'd386: inv_x_count_next = 16'b0000000010101010; // 1/386 = 0.0025906736
//      10'd387: inv_x_count_next = 16'b0000000010101001; // 1/387 = 0.0025839793
//      10'd388: inv_x_count_next = 16'b0000000010101001; // 1/388 = 0.0025773196
//      10'd389: inv_x_count_next = 16'b0000000010101000; // 1/389 = 0.0025706941
//      10'd390: inv_x_count_next = 16'b0000000010101000; // 1/390 = 0.0025641026
//      10'd391: inv_x_count_next = 16'b0000000010101000; // 1/391 = 0.0025575448
//      10'd392: inv_x_count_next = 16'b0000000010100111; // 1/392 = 0.0025510204
//      10'd393: inv_x_count_next = 16'b0000000010100111; // 1/393 = 0.0025445293
//      10'd394: inv_x_count_next = 16'b0000000010100110; // 1/394 = 0.0025380711
//      10'd395: inv_x_count_next = 16'b0000000010100110; // 1/395 = 0.0025316456
//      10'd396: inv_x_count_next = 16'b0000000010100101; // 1/396 = 0.0025252525
//      10'd397: inv_x_count_next = 16'b0000000010100101; // 1/397 = 0.0025188917
//      10'd398: inv_x_count_next = 16'b0000000010100101; // 1/398 = 0.0025125628
//      10'd399: inv_x_count_next = 16'b0000000010100100; // 1/399 = 0.0025062657
//      10'd400: inv_x_count_next = 16'b0000000010100100; // 1/400 = 0.0025000000
//      10'd401: inv_x_count_next = 16'b0000000010100011; // 1/401 = 0.0024937656
//      10'd402: inv_x_count_next = 16'b0000000010100011; // 1/402 = 0.0024875622
//      10'd403: inv_x_count_next = 16'b0000000010100011; // 1/403 = 0.0024813896
//      10'd404: inv_x_count_next = 16'b0000000010100010; // 1/404 = 0.0024752475
//      10'd405: inv_x_count_next = 16'b0000000010100010; // 1/405 = 0.0024691358
//      10'd406: inv_x_count_next = 16'b0000000010100001; // 1/406 = 0.0024630542
//      10'd407: inv_x_count_next = 16'b0000000010100001; // 1/407 = 0.0024570025
//      10'd408: inv_x_count_next = 16'b0000000010100001; // 1/408 = 0.0024509804
//      10'd409: inv_x_count_next = 16'b0000000010100000; // 1/409 = 0.0024449878
//      10'd410: inv_x_count_next = 16'b0000000010100000; // 1/410 = 0.0024390244
//      10'd411: inv_x_count_next = 16'b0000000010011111; // 1/411 = 0.0024330900
//      10'd412: inv_x_count_next = 16'b0000000010011111; // 1/412 = 0.0024271845
//      10'd413: inv_x_count_next = 16'b0000000010011111; // 1/413 = 0.0024213075
//      10'd414: inv_x_count_next = 16'b0000000010011110; // 1/414 = 0.0024154589
//      10'd415: inv_x_count_next = 16'b0000000010011110; // 1/415 = 0.0024096386
//      10'd416: inv_x_count_next = 16'b0000000010011110; // 1/416 = 0.0024038462
//      10'd417: inv_x_count_next = 16'b0000000010011101; // 1/417 = 0.0023980815
//      10'd418: inv_x_count_next = 16'b0000000010011101; // 1/418 = 0.0023923445
//      10'd419: inv_x_count_next = 16'b0000000010011100; // 1/419 = 0.0023866348
//      10'd420: inv_x_count_next = 16'b0000000010011100; // 1/420 = 0.0023809524
//      10'd421: inv_x_count_next = 16'b0000000010011100; // 1/421 = 0.0023752969
//      10'd422: inv_x_count_next = 16'b0000000010011011; // 1/422 = 0.0023696682
//      10'd423: inv_x_count_next = 16'b0000000010011011; // 1/423 = 0.0023640662
//      10'd424: inv_x_count_next = 16'b0000000010011011; // 1/424 = 0.0023584906
//      10'd425: inv_x_count_next = 16'b0000000010011010; // 1/425 = 0.0023529412
//      10'd426: inv_x_count_next = 16'b0000000010011010; // 1/426 = 0.0023474178
//      10'd427: inv_x_count_next = 16'b0000000010011001; // 1/427 = 0.0023419204
//      10'd428: inv_x_count_next = 16'b0000000010011001; // 1/428 = 0.0023364486
//      10'd429: inv_x_count_next = 16'b0000000010011001; // 1/429 = 0.0023310023
//      10'd430: inv_x_count_next = 16'b0000000010011000; // 1/430 = 0.0023255814
//      10'd431: inv_x_count_next = 16'b0000000010011000; // 1/431 = 0.0023201856
//      10'd432: inv_x_count_next = 16'b0000000010011000; // 1/432 = 0.0023148148
//      10'd433: inv_x_count_next = 16'b0000000010010111; // 1/433 = 0.0023094688
//      10'd434: inv_x_count_next = 16'b0000000010010111; // 1/434 = 0.0023041475
//      10'd435: inv_x_count_next = 16'b0000000010010111; // 1/435 = 0.0022988506
//      10'd436: inv_x_count_next = 16'b0000000010010110; // 1/436 = 0.0022935780
//      10'd437: inv_x_count_next = 16'b0000000010010110; // 1/437 = 0.0022883295
//      10'd438: inv_x_count_next = 16'b0000000010010110; // 1/438 = 0.0022831050
//      10'd439: inv_x_count_next = 16'b0000000010010101; // 1/439 = 0.0022779043
//      10'd440: inv_x_count_next = 16'b0000000010010101; // 1/440 = 0.0022727273
//      10'd441: inv_x_count_next = 16'b0000000010010101; // 1/441 = 0.0022675737
//      10'd442: inv_x_count_next = 16'b0000000010010100; // 1/442 = 0.0022624434
//      10'd443: inv_x_count_next = 16'b0000000010010100; // 1/443 = 0.0022573363
//      10'd444: inv_x_count_next = 16'b0000000010010100; // 1/444 = 0.0022522523
//      10'd445: inv_x_count_next = 16'b0000000010010011; // 1/445 = 0.0022471910
//      10'd446: inv_x_count_next = 16'b0000000010010011; // 1/446 = 0.0022421525
//      10'd447: inv_x_count_next = 16'b0000000010010011; // 1/447 = 0.0022371365
//      10'd448: inv_x_count_next = 16'b0000000010010010; // 1/448 = 0.0022321429
//      10'd449: inv_x_count_next = 16'b0000000010010010; // 1/449 = 0.0022271715
//      10'd450: inv_x_count_next = 16'b0000000010010010; // 1/450 = 0.0022222222
//      10'd451: inv_x_count_next = 16'b0000000010010001; // 1/451 = 0.0022172949
//      10'd452: inv_x_count_next = 16'b0000000010010001; // 1/452 = 0.0022123894
//      10'd453: inv_x_count_next = 16'b0000000010010001; // 1/453 = 0.0022075055
//      10'd454: inv_x_count_next = 16'b0000000010010000; // 1/454 = 0.0022026432
//      10'd455: inv_x_count_next = 16'b0000000010010000; // 1/455 = 0.0021978022
//      10'd456: inv_x_count_next = 16'b0000000010010000; // 1/456 = 0.0021929825
//      10'd457: inv_x_count_next = 16'b0000000010001111; // 1/457 = 0.0021881838
//      10'd458: inv_x_count_next = 16'b0000000010001111; // 1/458 = 0.0021834061
//      10'd459: inv_x_count_next = 16'b0000000010001111; // 1/459 = 0.0021786492
//      10'd460: inv_x_count_next = 16'b0000000010001110; // 1/460 = 0.0021739130
//      10'd461: inv_x_count_next = 16'b0000000010001110; // 1/461 = 0.0021691974
//      10'd462: inv_x_count_next = 16'b0000000010001110; // 1/462 = 0.0021645022
//      10'd463: inv_x_count_next = 16'b0000000010001110; // 1/463 = 0.0021598272
//      10'd464: inv_x_count_next = 16'b0000000010001101; // 1/464 = 0.0021551724
//      10'd465: inv_x_count_next = 16'b0000000010001101; // 1/465 = 0.0021505376
//      10'd466: inv_x_count_next = 16'b0000000010001101; // 1/466 = 0.0021459227
//      10'd467: inv_x_count_next = 16'b0000000010001100; // 1/467 = 0.0021413276
//      10'd468: inv_x_count_next = 16'b0000000010001100; // 1/468 = 0.0021367521
//      10'd469: inv_x_count_next = 16'b0000000010001100; // 1/469 = 0.0021321962
//      10'd470: inv_x_count_next = 16'b0000000010001011; // 1/470 = 0.0021276596
//      10'd471: inv_x_count_next = 16'b0000000010001011; // 1/471 = 0.0021231423
//      10'd472: inv_x_count_next = 16'b0000000010001011; // 1/472 = 0.0021186441
//      10'd473: inv_x_count_next = 16'b0000000010001011; // 1/473 = 0.0021141649
//      10'd474: inv_x_count_next = 16'b0000000010001010; // 1/474 = 0.0021097046
//      10'd475: inv_x_count_next = 16'b0000000010001010; // 1/475 = 0.0021052632
//      10'd476: inv_x_count_next = 16'b0000000010001010; // 1/476 = 0.0021008403
//      10'd477: inv_x_count_next = 16'b0000000010001001; // 1/477 = 0.0020964361
//      10'd478: inv_x_count_next = 16'b0000000010001001; // 1/478 = 0.0020920502
//      10'd479: inv_x_count_next = 16'b0000000010001001; // 1/479 = 0.0020876827
//      10'd480: inv_x_count_next = 16'b0000000010001001; // 1/480 = 0.0020833333
//      10'd481: inv_x_count_next = 16'b0000000010001000; // 1/481 = 0.0020790021
//      10'd482: inv_x_count_next = 16'b0000000010001000; // 1/482 = 0.0020746888
//      10'd483: inv_x_count_next = 16'b0000000010001000; // 1/483 = 0.0020703934
//      10'd484: inv_x_count_next = 16'b0000000010000111; // 1/484 = 0.0020661157
//      10'd485: inv_x_count_next = 16'b0000000010000111; // 1/485 = 0.0020618557
//      10'd486: inv_x_count_next = 16'b0000000010000111; // 1/486 = 0.0020576132
//      10'd487: inv_x_count_next = 16'b0000000010000111; // 1/487 = 0.0020533881
//      10'd488: inv_x_count_next = 16'b0000000010000110; // 1/488 = 0.0020491803
//      10'd489: inv_x_count_next = 16'b0000000010000110; // 1/489 = 0.0020449898
//      10'd490: inv_x_count_next = 16'b0000000010000110; // 1/490 = 0.0020408163
//      10'd491: inv_x_count_next = 16'b0000000010000101; // 1/491 = 0.0020366599
//      10'd492: inv_x_count_next = 16'b0000000010000101; // 1/492 = 0.0020325203
//      10'd493: inv_x_count_next = 16'b0000000010000101; // 1/493 = 0.0020283976
//      10'd494: inv_x_count_next = 16'b0000000010000101; // 1/494 = 0.0020242915
//      10'd495: inv_x_count_next = 16'b0000000010000100; // 1/495 = 0.0020202020
//      10'd496: inv_x_count_next = 16'b0000000010000100; // 1/496 = 0.0020161290
//      10'd497: inv_x_count_next = 16'b0000000010000100; // 1/497 = 0.0020120724
//      10'd498: inv_x_count_next = 16'b0000000010000100; // 1/498 = 0.0020080321
//      10'd499: inv_x_count_next = 16'b0000000010000011; // 1/499 = 0.0020040080
//      10'd500: inv_x_count_next = 16'b0000000010000011; // 1/500 = 0.0020000000
//      10'd501: inv_x_count_next = 16'b0000000010000011; // 1/501 = 0.0019960080
//      10'd502: inv_x_count_next = 16'b0000000010000011; // 1/502 = 0.0019920319
//      10'd503: inv_x_count_next = 16'b0000000010000010; // 1/503 = 0.0019880716
//      10'd504: inv_x_count_next = 16'b0000000010000010; // 1/504 = 0.0019841270
//      10'd505: inv_x_count_next = 16'b0000000010000010; // 1/505 = 0.0019801980
//      10'd506: inv_x_count_next = 16'b0000000010000010; // 1/506 = 0.0019762846
//      10'd507: inv_x_count_next = 16'b0000000010000001; // 1/507 = 0.0019723866
//      10'd508: inv_x_count_next = 16'b0000000010000001; // 1/508 = 0.0019685039
//      10'd509: inv_x_count_next = 16'b0000000010000001; // 1/509 = 0.0019646365
//      10'd510: inv_x_count_next = 16'b0000000010000001; // 1/510 = 0.0019607843
//      10'd511: inv_x_count_next = 16'b0000000010000000; // 1/511 = 0.0019569472
//      10'd512: inv_x_count_next = 16'b0000000010000000; // 1/512 = 0.0019531250
//      10'd513: inv_x_count_next = 16'b0000000010000000; // 1/513 = 0.0019493177
//      10'd514: inv_x_count_next = 16'b0000000010000000; // 1/514 = 0.0019455253
//      10'd515: inv_x_count_next = 16'b0000000001111111; // 1/515 = 0.0019417476
//      10'd516: inv_x_count_next = 16'b0000000001111111; // 1/516 = 0.0019379845
//      10'd517: inv_x_count_next = 16'b0000000001111111; // 1/517 = 0.0019342360
//      10'd518: inv_x_count_next = 16'b0000000001111111; // 1/518 = 0.0019305019
//      10'd519: inv_x_count_next = 16'b0000000001111110; // 1/519 = 0.0019267823
//      10'd520: inv_x_count_next = 16'b0000000001111110; // 1/520 = 0.0019230769
//      10'd521: inv_x_count_next = 16'b0000000001111110; // 1/521 = 0.0019193858
//      10'd522: inv_x_count_next = 16'b0000000001111110; // 1/522 = 0.0019157088
//      10'd523: inv_x_count_next = 16'b0000000001111101; // 1/523 = 0.0019120459
//      10'd524: inv_x_count_next = 16'b0000000001111101; // 1/524 = 0.0019083969
//      10'd525: inv_x_count_next = 16'b0000000001111101; // 1/525 = 0.0019047619
//      10'd526: inv_x_count_next = 16'b0000000001111101; // 1/526 = 0.0019011407
//      10'd527: inv_x_count_next = 16'b0000000001111100; // 1/527 = 0.0018975332
//      10'd528: inv_x_count_next = 16'b0000000001111100; // 1/528 = 0.0018939394
//      10'd529: inv_x_count_next = 16'b0000000001111100; // 1/529 = 0.0018903592
//      10'd530: inv_x_count_next = 16'b0000000001111100; // 1/530 = 0.0018867925
//      10'd531: inv_x_count_next = 16'b0000000001111011; // 1/531 = 0.0018832392
//      10'd532: inv_x_count_next = 16'b0000000001111011; // 1/532 = 0.0018796992
//      10'd533: inv_x_count_next = 16'b0000000001111011; // 1/533 = 0.0018761726
//      10'd534: inv_x_count_next = 16'b0000000001111011; // 1/534 = 0.0018726592
//      10'd535: inv_x_count_next = 16'b0000000001111010; // 1/535 = 0.0018691589
//      10'd536: inv_x_count_next = 16'b0000000001111010; // 1/536 = 0.0018656716
//      10'd537: inv_x_count_next = 16'b0000000001111010; // 1/537 = 0.0018621974
//      10'd538: inv_x_count_next = 16'b0000000001111010; // 1/538 = 0.0018587361
//      10'd539: inv_x_count_next = 16'b0000000001111010; // 1/539 = 0.0018552876
//      10'd540: inv_x_count_next = 16'b0000000001111001; // 1/540 = 0.0018518519
//      10'd541: inv_x_count_next = 16'b0000000001111001; // 1/541 = 0.0018484288
//      10'd542: inv_x_count_next = 16'b0000000001111001; // 1/542 = 0.0018450185
//      10'd543: inv_x_count_next = 16'b0000000001111001; // 1/543 = 0.0018416206
//      10'd544: inv_x_count_next = 16'b0000000001111000; // 1/544 = 0.0018382353
//      10'd545: inv_x_count_next = 16'b0000000001111000; // 1/545 = 0.0018348624
//      10'd546: inv_x_count_next = 16'b0000000001111000; // 1/546 = 0.0018315018
//      10'd547: inv_x_count_next = 16'b0000000001111000; // 1/547 = 0.0018281536
//      10'd548: inv_x_count_next = 16'b0000000001111000; // 1/548 = 0.0018248175
//      10'd549: inv_x_count_next = 16'b0000000001110111; // 1/549 = 0.0018214936
//      10'd550: inv_x_count_next = 16'b0000000001110111; // 1/550 = 0.0018181818
//      10'd551: inv_x_count_next = 16'b0000000001110111; // 1/551 = 0.0018148820
//      10'd552: inv_x_count_next = 16'b0000000001110111; // 1/552 = 0.0018115942
//      10'd553: inv_x_count_next = 16'b0000000001110111; // 1/553 = 0.0018083183
//      10'd554: inv_x_count_next = 16'b0000000001110110; // 1/554 = 0.0018050542
//      10'd555: inv_x_count_next = 16'b0000000001110110; // 1/555 = 0.0018018018
//      10'd556: inv_x_count_next = 16'b0000000001110110; // 1/556 = 0.0017985612
//      10'd557: inv_x_count_next = 16'b0000000001110110; // 1/557 = 0.0017953321
//      10'd558: inv_x_count_next = 16'b0000000001110101; // 1/558 = 0.0017921147
//      10'd559: inv_x_count_next = 16'b0000000001110101; // 1/559 = 0.0017889088
//      10'd560: inv_x_count_next = 16'b0000000001110101; // 1/560 = 0.0017857143
//      10'd561: inv_x_count_next = 16'b0000000001110101; // 1/561 = 0.0017825312
//      10'd562: inv_x_count_next = 16'b0000000001110101; // 1/562 = 0.0017793594
//      10'd563: inv_x_count_next = 16'b0000000001110100; // 1/563 = 0.0017761989
//      10'd564: inv_x_count_next = 16'b0000000001110100; // 1/564 = 0.0017730496
//      10'd565: inv_x_count_next = 16'b0000000001110100; // 1/565 = 0.0017699115
//      10'd566: inv_x_count_next = 16'b0000000001110100; // 1/566 = 0.0017667845
//      10'd567: inv_x_count_next = 16'b0000000001110100; // 1/567 = 0.0017636684
//      10'd568: inv_x_count_next = 16'b0000000001110011; // 1/568 = 0.0017605634
//      10'd569: inv_x_count_next = 16'b0000000001110011; // 1/569 = 0.0017574692
//      10'd570: inv_x_count_next = 16'b0000000001110011; // 1/570 = 0.0017543860
//      10'd571: inv_x_count_next = 16'b0000000001110011; // 1/571 = 0.0017513135
//      10'd572: inv_x_count_next = 16'b0000000001110011; // 1/572 = 0.0017482517
//      10'd573: inv_x_count_next = 16'b0000000001110010; // 1/573 = 0.0017452007
//      10'd574: inv_x_count_next = 16'b0000000001110010; // 1/574 = 0.0017421603
//      10'd575: inv_x_count_next = 16'b0000000001110010; // 1/575 = 0.0017391304
//      10'd576: inv_x_count_next = 16'b0000000001110010; // 1/576 = 0.0017361111
//      10'd577: inv_x_count_next = 16'b0000000001110010; // 1/577 = 0.0017331023
//      10'd578: inv_x_count_next = 16'b0000000001110001; // 1/578 = 0.0017301038
//      10'd579: inv_x_count_next = 16'b0000000001110001; // 1/579 = 0.0017271157
//      10'd580: inv_x_count_next = 16'b0000000001110001; // 1/580 = 0.0017241379
//      10'd581: inv_x_count_next = 16'b0000000001110001; // 1/581 = 0.0017211704
//      10'd582: inv_x_count_next = 16'b0000000001110001; // 1/582 = 0.0017182131
//      10'd583: inv_x_count_next = 16'b0000000001110000; // 1/583 = 0.0017152659
//      10'd584: inv_x_count_next = 16'b0000000001110000; // 1/584 = 0.0017123288
//      10'd585: inv_x_count_next = 16'b0000000001110000; // 1/585 = 0.0017094017
//      10'd586: inv_x_count_next = 16'b0000000001110000; // 1/586 = 0.0017064846
//      10'd587: inv_x_count_next = 16'b0000000001110000; // 1/587 = 0.0017035775
//      10'd588: inv_x_count_next = 16'b0000000001101111; // 1/588 = 0.0017006803
//      10'd589: inv_x_count_next = 16'b0000000001101111; // 1/589 = 0.0016977929
//      10'd590: inv_x_count_next = 16'b0000000001101111; // 1/590 = 0.0016949153
//      10'd591: inv_x_count_next = 16'b0000000001101111; // 1/591 = 0.0016920474
//      10'd592: inv_x_count_next = 16'b0000000001101111; // 1/592 = 0.0016891892
//      10'd593: inv_x_count_next = 16'b0000000001101111; // 1/593 = 0.0016863406
//      10'd594: inv_x_count_next = 16'b0000000001101110; // 1/594 = 0.0016835017
//      10'd595: inv_x_count_next = 16'b0000000001101110; // 1/595 = 0.0016806723
//      10'd596: inv_x_count_next = 16'b0000000001101110; // 1/596 = 0.0016778523
//      10'd597: inv_x_count_next = 16'b0000000001101110; // 1/597 = 0.0016750419
//      10'd598: inv_x_count_next = 16'b0000000001101110; // 1/598 = 0.0016722408
//      10'd599: inv_x_count_next = 16'b0000000001101101; // 1/599 = 0.0016694491
//      10'd600: inv_x_count_next = 16'b0000000001101101; // 1/600 = 0.0016666667
//      10'd601: inv_x_count_next = 16'b0000000001101101; // 1/601 = 0.0016638935
//      10'd602: inv_x_count_next = 16'b0000000001101101; // 1/602 = 0.0016611296
//      10'd603: inv_x_count_next = 16'b0000000001101101; // 1/603 = 0.0016583748
//      10'd604: inv_x_count_next = 16'b0000000001101101; // 1/604 = 0.0016556291
//      10'd605: inv_x_count_next = 16'b0000000001101100; // 1/605 = 0.0016528926
//      10'd606: inv_x_count_next = 16'b0000000001101100; // 1/606 = 0.0016501650
//      10'd607: inv_x_count_next = 16'b0000000001101100; // 1/607 = 0.0016474465
//      10'd608: inv_x_count_next = 16'b0000000001101100; // 1/608 = 0.0016447368
//      10'd609: inv_x_count_next = 16'b0000000001101100; // 1/609 = 0.0016420361
//      10'd610: inv_x_count_next = 16'b0000000001101011; // 1/610 = 0.0016393443
//      10'd611: inv_x_count_next = 16'b0000000001101011; // 1/611 = 0.0016366612
//      10'd612: inv_x_count_next = 16'b0000000001101011; // 1/612 = 0.0016339869
//      10'd613: inv_x_count_next = 16'b0000000001101011; // 1/613 = 0.0016313214
//      10'd614: inv_x_count_next = 16'b0000000001101011; // 1/614 = 0.0016286645
//      10'd615: inv_x_count_next = 16'b0000000001101011; // 1/615 = 0.0016260163
//      10'd616: inv_x_count_next = 16'b0000000001101010; // 1/616 = 0.0016233766
//      10'd617: inv_x_count_next = 16'b0000000001101010; // 1/617 = 0.0016207455
//      10'd618: inv_x_count_next = 16'b0000000001101010; // 1/618 = 0.0016181230
//      10'd619: inv_x_count_next = 16'b0000000001101010; // 1/619 = 0.0016155089
//      10'd620: inv_x_count_next = 16'b0000000001101010; // 1/620 = 0.0016129032
//      10'd621: inv_x_count_next = 16'b0000000001101010; // 1/621 = 0.0016103060
//      10'd622: inv_x_count_next = 16'b0000000001101001; // 1/622 = 0.0016077170
//      10'd623: inv_x_count_next = 16'b0000000001101001; // 1/623 = 0.0016051364
//      10'd624: inv_x_count_next = 16'b0000000001101001; // 1/624 = 0.0016025641
//      10'd625: inv_x_count_next = 16'b0000000001101001; // 1/625 = 0.0016000000
//      10'd626: inv_x_count_next = 16'b0000000001101001; // 1/626 = 0.0015974441
//      10'd627: inv_x_count_next = 16'b0000000001101001; // 1/627 = 0.0015948963
//      10'd628: inv_x_count_next = 16'b0000000001101000; // 1/628 = 0.0015923567
//      10'd629: inv_x_count_next = 16'b0000000001101000; // 1/629 = 0.0015898251
//      10'd630: inv_x_count_next = 16'b0000000001101000; // 1/630 = 0.0015873016
//      10'd631: inv_x_count_next = 16'b0000000001101000; // 1/631 = 0.0015847861
//      10'd632: inv_x_count_next = 16'b0000000001101000; // 1/632 = 0.0015822785
//      10'd633: inv_x_count_next = 16'b0000000001101000; // 1/633 = 0.0015797788
//      10'd634: inv_x_count_next = 16'b0000000001100111; // 1/634 = 0.0015772871
//      10'd635: inv_x_count_next = 16'b0000000001100111; // 1/635 = 0.0015748031
//      10'd636: inv_x_count_next = 16'b0000000001100111; // 1/636 = 0.0015723270
//      10'd637: inv_x_count_next = 16'b0000000001100111; // 1/637 = 0.0015698587
//      10'd638: inv_x_count_next = 16'b0000000001100111; // 1/638 = 0.0015673981
//      10'd639: inv_x_count_next = 16'b0000000001100111; // 1/639 = 0.0015649452
//      10'd640: inv_x_count_next = 16'b0000000001100110; // 1/640 = 0.0015625000
//      10'd641: inv_x_count_next = 16'b0000000001100110; // 1/641 = 0.0015600624
//      10'd642: inv_x_count_next = 16'b0000000001100110; // 1/642 = 0.0015576324
//      10'd643: inv_x_count_next = 16'b0000000001100110; // 1/643 = 0.0015552100
//      10'd644: inv_x_count_next = 16'b0000000001100110; // 1/644 = 0.0015527950
//      10'd645: inv_x_count_next = 16'b0000000001100110; // 1/645 = 0.0015503876
//      10'd646: inv_x_count_next = 16'b0000000001100101; // 1/646 = 0.0015479876
//      10'd647: inv_x_count_next = 16'b0000000001100101; // 1/647 = 0.0015455951
//      10'd648: inv_x_count_next = 16'b0000000001100101; // 1/648 = 0.0015432099
//      10'd649: inv_x_count_next = 16'b0000000001100101; // 1/649 = 0.0015408320
//      10'd650: inv_x_count_next = 16'b0000000001100101; // 1/650 = 0.0015384615
//      10'd651: inv_x_count_next = 16'b0000000001100101; // 1/651 = 0.0015360983
//      10'd652: inv_x_count_next = 16'b0000000001100101; // 1/652 = 0.0015337423
//      10'd653: inv_x_count_next = 16'b0000000001100100; // 1/653 = 0.0015313936
//      10'd654: inv_x_count_next = 16'b0000000001100100; // 1/654 = 0.0015290520
//      10'd655: inv_x_count_next = 16'b0000000001100100; // 1/655 = 0.0015267176
//      10'd656: inv_x_count_next = 16'b0000000001100100; // 1/656 = 0.0015243902
//      10'd657: inv_x_count_next = 16'b0000000001100100; // 1/657 = 0.0015220700
//      10'd658: inv_x_count_next = 16'b0000000001100100; // 1/658 = 0.0015197568
//      10'd659: inv_x_count_next = 16'b0000000001100011; // 1/659 = 0.0015174507
//      10'd660: inv_x_count_next = 16'b0000000001100011; // 1/660 = 0.0015151515
//      10'd661: inv_x_count_next = 16'b0000000001100011; // 1/661 = 0.0015128593
//      10'd662: inv_x_count_next = 16'b0000000001100011; // 1/662 = 0.0015105740
//      10'd663: inv_x_count_next = 16'b0000000001100011; // 1/663 = 0.0015082956
//      10'd664: inv_x_count_next = 16'b0000000001100011; // 1/664 = 0.0015060241
//      10'd665: inv_x_count_next = 16'b0000000001100011; // 1/665 = 0.0015037594
//      10'd666: inv_x_count_next = 16'b0000000001100010; // 1/666 = 0.0015015015
//      10'd667: inv_x_count_next = 16'b0000000001100010; // 1/667 = 0.0014992504
//      10'd668: inv_x_count_next = 16'b0000000001100010; // 1/668 = 0.0014970060
//      10'd669: inv_x_count_next = 16'b0000000001100010; // 1/669 = 0.0014947683
//      10'd670: inv_x_count_next = 16'b0000000001100010; // 1/670 = 0.0014925373
//      10'd671: inv_x_count_next = 16'b0000000001100010; // 1/671 = 0.0014903130
//      10'd672: inv_x_count_next = 16'b0000000001100010; // 1/672 = 0.0014880952
//      10'd673: inv_x_count_next = 16'b0000000001100001; // 1/673 = 0.0014858841
//      10'd674: inv_x_count_next = 16'b0000000001100001; // 1/674 = 0.0014836795
//      10'd675: inv_x_count_next = 16'b0000000001100001; // 1/675 = 0.0014814815
//      10'd676: inv_x_count_next = 16'b0000000001100001; // 1/676 = 0.0014792899
//      10'd677: inv_x_count_next = 16'b0000000001100001; // 1/677 = 0.0014771049
//      10'd678: inv_x_count_next = 16'b0000000001100001; // 1/678 = 0.0014749263
//      10'd679: inv_x_count_next = 16'b0000000001100001; // 1/679 = 0.0014727541
//      10'd680: inv_x_count_next = 16'b0000000001100000; // 1/680 = 0.0014705882
//      10'd681: inv_x_count_next = 16'b0000000001100000; // 1/681 = 0.0014684288
//      10'd682: inv_x_count_next = 16'b0000000001100000; // 1/682 = 0.0014662757
//      10'd683: inv_x_count_next = 16'b0000000001100000; // 1/683 = 0.0014641288
//      10'd684: inv_x_count_next = 16'b0000000001100000; // 1/684 = 0.0014619883
//      10'd685: inv_x_count_next = 16'b0000000001100000; // 1/685 = 0.0014598540
//      10'd686: inv_x_count_next = 16'b0000000001100000; // 1/686 = 0.0014577259
//      10'd687: inv_x_count_next = 16'b0000000001011111; // 1/687 = 0.0014556041
//      10'd688: inv_x_count_next = 16'b0000000001011111; // 1/688 = 0.0014534884
//      10'd689: inv_x_count_next = 16'b0000000001011111; // 1/689 = 0.0014513788
//      10'd690: inv_x_count_next = 16'b0000000001011111; // 1/690 = 0.0014492754
//      10'd691: inv_x_count_next = 16'b0000000001011111; // 1/691 = 0.0014471780
//      10'd692: inv_x_count_next = 16'b0000000001011111; // 1/692 = 0.0014450867
//      10'd693: inv_x_count_next = 16'b0000000001011111; // 1/693 = 0.0014430014
//      10'd694: inv_x_count_next = 16'b0000000001011110; // 1/694 = 0.0014409222
//      10'd695: inv_x_count_next = 16'b0000000001011110; // 1/695 = 0.0014388489
//      10'd696: inv_x_count_next = 16'b0000000001011110; // 1/696 = 0.0014367816
//      10'd697: inv_x_count_next = 16'b0000000001011110; // 1/697 = 0.0014347202
//      10'd698: inv_x_count_next = 16'b0000000001011110; // 1/698 = 0.0014326648
//      10'd699: inv_x_count_next = 16'b0000000001011110; // 1/699 = 0.0014306152
//      10'd700: inv_x_count_next = 16'b0000000001011110; // 1/700 = 0.0014285714
//      10'd701: inv_x_count_next = 16'b0000000001011101; // 1/701 = 0.0014265335
//      10'd702: inv_x_count_next = 16'b0000000001011101; // 1/702 = 0.0014245014
//      10'd703: inv_x_count_next = 16'b0000000001011101; // 1/703 = 0.0014224751
//      10'd704: inv_x_count_next = 16'b0000000001011101; // 1/704 = 0.0014204545
//      10'd705: inv_x_count_next = 16'b0000000001011101; // 1/705 = 0.0014184397
//      10'd706: inv_x_count_next = 16'b0000000001011101; // 1/706 = 0.0014164306
//      10'd707: inv_x_count_next = 16'b0000000001011101; // 1/707 = 0.0014144272
//      10'd708: inv_x_count_next = 16'b0000000001011101; // 1/708 = 0.0014124294
//      10'd709: inv_x_count_next = 16'b0000000001011100; // 1/709 = 0.0014104372
//      10'd710: inv_x_count_next = 16'b0000000001011100; // 1/710 = 0.0014084507
//      10'd711: inv_x_count_next = 16'b0000000001011100; // 1/711 = 0.0014064698
//      10'd712: inv_x_count_next = 16'b0000000001011100; // 1/712 = 0.0014044944
//      10'd713: inv_x_count_next = 16'b0000000001011100; // 1/713 = 0.0014025245
//      10'd714: inv_x_count_next = 16'b0000000001011100; // 1/714 = 0.0014005602
//      10'd715: inv_x_count_next = 16'b0000000001011100; // 1/715 = 0.0013986014
//      10'd716: inv_x_count_next = 16'b0000000001011100; // 1/716 = 0.0013966480
//      10'd717: inv_x_count_next = 16'b0000000001011011; // 1/717 = 0.0013947001
//      10'd718: inv_x_count_next = 16'b0000000001011011; // 1/718 = 0.0013927577
//      10'd719: inv_x_count_next = 16'b0000000001011011; // 1/719 = 0.0013908206
//      10'd720: inv_x_count_next = 16'b0000000001011011; // 1/720 = 0.0013888889
//      10'd721: inv_x_count_next = 16'b0000000001011011; // 1/721 = 0.0013869626
//      10'd722: inv_x_count_next = 16'b0000000001011011; // 1/722 = 0.0013850416
//      10'd723: inv_x_count_next = 16'b0000000001011011; // 1/723 = 0.0013831259
//      10'd724: inv_x_count_next = 16'b0000000001011011; // 1/724 = 0.0013812155
//      10'd725: inv_x_count_next = 16'b0000000001011010; // 1/725 = 0.0013793103
//      10'd726: inv_x_count_next = 16'b0000000001011010; // 1/726 = 0.0013774105
//      10'd727: inv_x_count_next = 16'b0000000001011010; // 1/727 = 0.0013755158
//      10'd728: inv_x_count_next = 16'b0000000001011010; // 1/728 = 0.0013736264
//      10'd729: inv_x_count_next = 16'b0000000001011010; // 1/729 = 0.0013717421
//      10'd730: inv_x_count_next = 16'b0000000001011010; // 1/730 = 0.0013698630
//      10'd731: inv_x_count_next = 16'b0000000001011010; // 1/731 = 0.0013679891
//      10'd732: inv_x_count_next = 16'b0000000001011010; // 1/732 = 0.0013661202
//      10'd733: inv_x_count_next = 16'b0000000001011001; // 1/733 = 0.0013642565
//      10'd734: inv_x_count_next = 16'b0000000001011001; // 1/734 = 0.0013623978
//      10'd735: inv_x_count_next = 16'b0000000001011001; // 1/735 = 0.0013605442
//      10'd736: inv_x_count_next = 16'b0000000001011001; // 1/736 = 0.0013586957
//      10'd737: inv_x_count_next = 16'b0000000001011001; // 1/737 = 0.0013568521
//      10'd738: inv_x_count_next = 16'b0000000001011001; // 1/738 = 0.0013550136
//      10'd739: inv_x_count_next = 16'b0000000001011001; // 1/739 = 0.0013531800
//      10'd740: inv_x_count_next = 16'b0000000001011001; // 1/740 = 0.0013513514
//      10'd741: inv_x_count_next = 16'b0000000001011000; // 1/741 = 0.0013495277
//      10'd742: inv_x_count_next = 16'b0000000001011000; // 1/742 = 0.0013477089
//      10'd743: inv_x_count_next = 16'b0000000001011000; // 1/743 = 0.0013458950
//      10'd744: inv_x_count_next = 16'b0000000001011000; // 1/744 = 0.0013440860
//      10'd745: inv_x_count_next = 16'b0000000001011000; // 1/745 = 0.0013422819
//      10'd746: inv_x_count_next = 16'b0000000001011000; // 1/746 = 0.0013404826
//      10'd747: inv_x_count_next = 16'b0000000001011000; // 1/747 = 0.0013386881
//      10'd748: inv_x_count_next = 16'b0000000001011000; // 1/748 = 0.0013368984
//      10'd749: inv_x_count_next = 16'b0000000001010111; // 1/749 = 0.0013351135
//      10'd750: inv_x_count_next = 16'b0000000001010111; // 1/750 = 0.0013333333
//      10'd751: inv_x_count_next = 16'b0000000001010111; // 1/751 = 0.0013315579
//      10'd752: inv_x_count_next = 16'b0000000001010111; // 1/752 = 0.0013297872
//      10'd753: inv_x_count_next = 16'b0000000001010111; // 1/753 = 0.0013280212
//      10'd754: inv_x_count_next = 16'b0000000001010111; // 1/754 = 0.0013262599
//      10'd755: inv_x_count_next = 16'b0000000001010111; // 1/755 = 0.0013245033
//      10'd756: inv_x_count_next = 16'b0000000001010111; // 1/756 = 0.0013227513
//      10'd757: inv_x_count_next = 16'b0000000001010111; // 1/757 = 0.0013210040
//      10'd758: inv_x_count_next = 16'b0000000001010110; // 1/758 = 0.0013192612
//      10'd759: inv_x_count_next = 16'b0000000001010110; // 1/759 = 0.0013175231
//      10'd760: inv_x_count_next = 16'b0000000001010110; // 1/760 = 0.0013157895
//      10'd761: inv_x_count_next = 16'b0000000001010110; // 1/761 = 0.0013140604
//      10'd762: inv_x_count_next = 16'b0000000001010110; // 1/762 = 0.0013123360
//      10'd763: inv_x_count_next = 16'b0000000001010110; // 1/763 = 0.0013106160
//      10'd764: inv_x_count_next = 16'b0000000001010110; // 1/764 = 0.0013089005
//      10'd765: inv_x_count_next = 16'b0000000001010110; // 1/765 = 0.0013071895
//      10'd766: inv_x_count_next = 16'b0000000001010110; // 1/766 = 0.0013054830
//      10'd767: inv_x_count_next = 16'b0000000001010101; // 1/767 = 0.0013037810
//      10'd768: inv_x_count_next = 16'b0000000001010101; // 1/768 = 0.0013020833
//      10'd769: inv_x_count_next = 16'b0000000001010101; // 1/769 = 0.0013003901
//      10'd770: inv_x_count_next = 16'b0000000001010101; // 1/770 = 0.0012987013
//      10'd771: inv_x_count_next = 16'b0000000001010101; // 1/771 = 0.0012970169
//      10'd772: inv_x_count_next = 16'b0000000001010101; // 1/772 = 0.0012953368
//      10'd773: inv_x_count_next = 16'b0000000001010101; // 1/773 = 0.0012936611
//      10'd774: inv_x_count_next = 16'b0000000001010101; // 1/774 = 0.0012919897
//      10'd775: inv_x_count_next = 16'b0000000001010101; // 1/775 = 0.0012903226
//      10'd776: inv_x_count_next = 16'b0000000001010100; // 1/776 = 0.0012886598
//      10'd777: inv_x_count_next = 16'b0000000001010100; // 1/777 = 0.0012870013
//      10'd778: inv_x_count_next = 16'b0000000001010100; // 1/778 = 0.0012853470
//      10'd779: inv_x_count_next = 16'b0000000001010100; // 1/779 = 0.0012836970
//      10'd780: inv_x_count_next = 16'b0000000001010100; // 1/780 = 0.0012820513
//      10'd781: inv_x_count_next = 16'b0000000001010100; // 1/781 = 0.0012804097
//      10'd782: inv_x_count_next = 16'b0000000001010100; // 1/782 = 0.0012787724
//      10'd783: inv_x_count_next = 16'b0000000001010100; // 1/783 = 0.0012771392
//      10'd784: inv_x_count_next = 16'b0000000001010100; // 1/784 = 0.0012755102
//      10'd785: inv_x_count_next = 16'b0000000001010011; // 1/785 = 0.0012738854
//      10'd786: inv_x_count_next = 16'b0000000001010011; // 1/786 = 0.0012722646
//      10'd787: inv_x_count_next = 16'b0000000001010011; // 1/787 = 0.0012706480
//      10'd788: inv_x_count_next = 16'b0000000001010011; // 1/788 = 0.0012690355
//      10'd789: inv_x_count_next = 16'b0000000001010011; // 1/789 = 0.0012674271
//      10'd790: inv_x_count_next = 16'b0000000001010011; // 1/790 = 0.0012658228
//      10'd791: inv_x_count_next = 16'b0000000001010011; // 1/791 = 0.0012642225
//      10'd792: inv_x_count_next = 16'b0000000001010011; // 1/792 = 0.0012626263
//      10'd793: inv_x_count_next = 16'b0000000001010011; // 1/793 = 0.0012610340
//      10'd794: inv_x_count_next = 16'b0000000001010011; // 1/794 = 0.0012594458
//      10'd795: inv_x_count_next = 16'b0000000001010010; // 1/795 = 0.0012578616
//      10'd796: inv_x_count_next = 16'b0000000001010010; // 1/796 = 0.0012562814
//      10'd797: inv_x_count_next = 16'b0000000001010010; // 1/797 = 0.0012547051
//      10'd798: inv_x_count_next = 16'b0000000001010010; // 1/798 = 0.0012531328
//      10'd799: inv_x_count_next = 16'b0000000001010010; // 1/799 = 0.0012515645
//      10'd800: inv_x_count_next = 16'b0000000001010010; // 1/800 = 0.0012500000
//      10'd801: inv_x_count_next = 16'b0000000001010010; // 1/801 = 0.0012484395
//      10'd802: inv_x_count_next = 16'b0000000001010010; // 1/802 = 0.0012468828
//      10'd803: inv_x_count_next = 16'b0000000001010010; // 1/803 = 0.0012453300
//      10'd804: inv_x_count_next = 16'b0000000001010010; // 1/804 = 0.0012437811
//      10'd805: inv_x_count_next = 16'b0000000001010001; // 1/805 = 0.0012422360
//      10'd806: inv_x_count_next = 16'b0000000001010001; // 1/806 = 0.0012406948
//      10'd807: inv_x_count_next = 16'b0000000001010001; // 1/807 = 0.0012391574
//      10'd808: inv_x_count_next = 16'b0000000001010001; // 1/808 = 0.0012376238
//      10'd809: inv_x_count_next = 16'b0000000001010001; // 1/809 = 0.0012360939
//      10'd810: inv_x_count_next = 16'b0000000001010001; // 1/810 = 0.0012345679
//      10'd811: inv_x_count_next = 16'b0000000001010001; // 1/811 = 0.0012330456
//      10'd812: inv_x_count_next = 16'b0000000001010001; // 1/812 = 0.0012315271
//      10'd813: inv_x_count_next = 16'b0000000001010001; // 1/813 = 0.0012300123
//      10'd814: inv_x_count_next = 16'b0000000001010001; // 1/814 = 0.0012285012
//      10'd815: inv_x_count_next = 16'b0000000001010000; // 1/815 = 0.0012269939
//      10'd816: inv_x_count_next = 16'b0000000001010000; // 1/816 = 0.0012254902
//      10'd817: inv_x_count_next = 16'b0000000001010000; // 1/817 = 0.0012239902
//      10'd818: inv_x_count_next = 16'b0000000001010000; // 1/818 = 0.0012224939
//      10'd819: inv_x_count_next = 16'b0000000001010000; // 1/819 = 0.0012210012
//      10'd820: inv_x_count_next = 16'b0000000001010000; // 1/820 = 0.0012195122
//      10'd821: inv_x_count_next = 16'b0000000001010000; // 1/821 = 0.0012180268
//      10'd822: inv_x_count_next = 16'b0000000001010000; // 1/822 = 0.0012165450
//      10'd823: inv_x_count_next = 16'b0000000001010000; // 1/823 = 0.0012150668
//      10'd824: inv_x_count_next = 16'b0000000001010000; // 1/824 = 0.0012135922
//      10'd825: inv_x_count_next = 16'b0000000001001111; // 1/825 = 0.0012121212
//      10'd826: inv_x_count_next = 16'b0000000001001111; // 1/826 = 0.0012106538
//      10'd827: inv_x_count_next = 16'b0000000001001111; // 1/827 = 0.0012091898
//      10'd828: inv_x_count_next = 16'b0000000001001111; // 1/828 = 0.0012077295
//      10'd829: inv_x_count_next = 16'b0000000001001111; // 1/829 = 0.0012062726
//      10'd830: inv_x_count_next = 16'b0000000001001111; // 1/830 = 0.0012048193
//      10'd831: inv_x_count_next = 16'b0000000001001111; // 1/831 = 0.0012033694
//      10'd832: inv_x_count_next = 16'b0000000001001111; // 1/832 = 0.0012019231
//      10'd833: inv_x_count_next = 16'b0000000001001111; // 1/833 = 0.0012004802
//      10'd834: inv_x_count_next = 16'b0000000001001111; // 1/834 = 0.0011990408
//      10'd835: inv_x_count_next = 16'b0000000001001110; // 1/835 = 0.0011976048
//      10'd836: inv_x_count_next = 16'b0000000001001110; // 1/836 = 0.0011961722
//      10'd837: inv_x_count_next = 16'b0000000001001110; // 1/837 = 0.0011947431
//      10'd838: inv_x_count_next = 16'b0000000001001110; // 1/838 = 0.0011933174
//      10'd839: inv_x_count_next = 16'b0000000001001110; // 1/839 = 0.0011918951
//      10'd840: inv_x_count_next = 16'b0000000001001110; // 1/840 = 0.0011904762
//      10'd841: inv_x_count_next = 16'b0000000001001110; // 1/841 = 0.0011890606
//      10'd842: inv_x_count_next = 16'b0000000001001110; // 1/842 = 0.0011876485
//      10'd843: inv_x_count_next = 16'b0000000001001110; // 1/843 = 0.0011862396
//      10'd844: inv_x_count_next = 16'b0000000001001110; // 1/844 = 0.0011848341
//      10'd845: inv_x_count_next = 16'b0000000001001110; // 1/845 = 0.0011834320
//      10'd846: inv_x_count_next = 16'b0000000001001101; // 1/846 = 0.0011820331
//      10'd847: inv_x_count_next = 16'b0000000001001101; // 1/847 = 0.0011806375
//      10'd848: inv_x_count_next = 16'b0000000001001101; // 1/848 = 0.0011792453
//      10'd849: inv_x_count_next = 16'b0000000001001101; // 1/849 = 0.0011778563
//      10'd850: inv_x_count_next = 16'b0000000001001101; // 1/850 = 0.0011764706
//      10'd851: inv_x_count_next = 16'b0000000001001101; // 1/851 = 0.0011750881
//      10'd852: inv_x_count_next = 16'b0000000001001101; // 1/852 = 0.0011737089
//      10'd853: inv_x_count_next = 16'b0000000001001101; // 1/853 = 0.0011723329
//      10'd854: inv_x_count_next = 16'b0000000001001101; // 1/854 = 0.0011709602
//      10'd855: inv_x_count_next = 16'b0000000001001101; // 1/855 = 0.0011695906
//      10'd856: inv_x_count_next = 16'b0000000001001101; // 1/856 = 0.0011682243
//      10'd857: inv_x_count_next = 16'b0000000001001100; // 1/857 = 0.0011668611
//      10'd858: inv_x_count_next = 16'b0000000001001100; // 1/858 = 0.0011655012
//      10'd859: inv_x_count_next = 16'b0000000001001100; // 1/859 = 0.0011641444
//      10'd860: inv_x_count_next = 16'b0000000001001100; // 1/860 = 0.0011627907
//      10'd861: inv_x_count_next = 16'b0000000001001100; // 1/861 = 0.0011614402
//      10'd862: inv_x_count_next = 16'b0000000001001100; // 1/862 = 0.0011600928
//      10'd863: inv_x_count_next = 16'b0000000001001100; // 1/863 = 0.0011587486
//      10'd864: inv_x_count_next = 16'b0000000001001100; // 1/864 = 0.0011574074
//      10'd865: inv_x_count_next = 16'b0000000001001100; // 1/865 = 0.0011560694
//      10'd866: inv_x_count_next = 16'b0000000001001100; // 1/866 = 0.0011547344
//      10'd867: inv_x_count_next = 16'b0000000001001100; // 1/867 = 0.0011534025
//      10'd868: inv_x_count_next = 16'b0000000001001100; // 1/868 = 0.0011520737
//      10'd869: inv_x_count_next = 16'b0000000001001011; // 1/869 = 0.0011507480
//      10'd870: inv_x_count_next = 16'b0000000001001011; // 1/870 = 0.0011494253
//      10'd871: inv_x_count_next = 16'b0000000001001011; // 1/871 = 0.0011481056
//      10'd872: inv_x_count_next = 16'b0000000001001011; // 1/872 = 0.0011467890
//      10'd873: inv_x_count_next = 16'b0000000001001011; // 1/873 = 0.0011454754
//      10'd874: inv_x_count_next = 16'b0000000001001011; // 1/874 = 0.0011441648
//      10'd875: inv_x_count_next = 16'b0000000001001011; // 1/875 = 0.0011428571
//      10'd876: inv_x_count_next = 16'b0000000001001011; // 1/876 = 0.0011415525
//      10'd877: inv_x_count_next = 16'b0000000001001011; // 1/877 = 0.0011402509
//      10'd878: inv_x_count_next = 16'b0000000001001011; // 1/878 = 0.0011389522
//      10'd879: inv_x_count_next = 16'b0000000001001011; // 1/879 = 0.0011376564
//      10'd880: inv_x_count_next = 16'b0000000001001010; // 1/880 = 0.0011363636
//      10'd881: inv_x_count_next = 16'b0000000001001010; // 1/881 = 0.0011350738
//      10'd882: inv_x_count_next = 16'b0000000001001010; // 1/882 = 0.0011337868
//      10'd883: inv_x_count_next = 16'b0000000001001010; // 1/883 = 0.0011325028
//      10'd884: inv_x_count_next = 16'b0000000001001010; // 1/884 = 0.0011312217
//      10'd885: inv_x_count_next = 16'b0000000001001010; // 1/885 = 0.0011299435
//      10'd886: inv_x_count_next = 16'b0000000001001010; // 1/886 = 0.0011286682
//      10'd887: inv_x_count_next = 16'b0000000001001010; // 1/887 = 0.0011273957
//      10'd888: inv_x_count_next = 16'b0000000001001010; // 1/888 = 0.0011261261
//      10'd889: inv_x_count_next = 16'b0000000001001010; // 1/889 = 0.0011248594
//      10'd890: inv_x_count_next = 16'b0000000001001010; // 1/890 = 0.0011235955
//      10'd891: inv_x_count_next = 16'b0000000001001010; // 1/891 = 0.0011223345
//      10'd892: inv_x_count_next = 16'b0000000001001001; // 1/892 = 0.0011210762
//      10'd893: inv_x_count_next = 16'b0000000001001001; // 1/893 = 0.0011198208
//      10'd894: inv_x_count_next = 16'b0000000001001001; // 1/894 = 0.0011185682
//      10'd895: inv_x_count_next = 16'b0000000001001001; // 1/895 = 0.0011173184
//      10'd896: inv_x_count_next = 16'b0000000001001001; // 1/896 = 0.0011160714
//      10'd897: inv_x_count_next = 16'b0000000001001001; // 1/897 = 0.0011148272
//      10'd898: inv_x_count_next = 16'b0000000001001001; // 1/898 = 0.0011135857
//      10'd899: inv_x_count_next = 16'b0000000001001001; // 1/899 = 0.0011123471
//      10'd900: inv_x_count_next = 16'b0000000001001001; // 1/900 = 0.0011111111
//      10'd901: inv_x_count_next = 16'b0000000001001001; // 1/901 = 0.0011098779
//      10'd902: inv_x_count_next = 16'b0000000001001001; // 1/902 = 0.0011086475
//      10'd903: inv_x_count_next = 16'b0000000001001001; // 1/903 = 0.0011074197
//      10'd904: inv_x_count_next = 16'b0000000001001000; // 1/904 = 0.0011061947
//      10'd905: inv_x_count_next = 16'b0000000001001000; // 1/905 = 0.0011049724
//      10'd906: inv_x_count_next = 16'b0000000001001000; // 1/906 = 0.0011037528
//      10'd907: inv_x_count_next = 16'b0000000001001000; // 1/907 = 0.0011025358
//      10'd908: inv_x_count_next = 16'b0000000001001000; // 1/908 = 0.0011013216
//      10'd909: inv_x_count_next = 16'b0000000001001000; // 1/909 = 0.0011001100
//      10'd910: inv_x_count_next = 16'b0000000001001000; // 1/910 = 0.0010989011
//      10'd911: inv_x_count_next = 16'b0000000001001000; // 1/911 = 0.0010976948
//      10'd912: inv_x_count_next = 16'b0000000001001000; // 1/912 = 0.0010964912
//      10'd913: inv_x_count_next = 16'b0000000001001000; // 1/913 = 0.0010952903
//      10'd914: inv_x_count_next = 16'b0000000001001000; // 1/914 = 0.0010940919
//      10'd915: inv_x_count_next = 16'b0000000001001000; // 1/915 = 0.0010928962
//      10'd916: inv_x_count_next = 16'b0000000001001000; // 1/916 = 0.0010917031
//      10'd917: inv_x_count_next = 16'b0000000001000111; // 1/917 = 0.0010905125
//      10'd918: inv_x_count_next = 16'b0000000001000111; // 1/918 = 0.0010893246
//      10'd919: inv_x_count_next = 16'b0000000001000111; // 1/919 = 0.0010881393
//      10'd920: inv_x_count_next = 16'b0000000001000111; // 1/920 = 0.0010869565
//      10'd921: inv_x_count_next = 16'b0000000001000111; // 1/921 = 0.0010857763
//      10'd922: inv_x_count_next = 16'b0000000001000111; // 1/922 = 0.0010845987
//      10'd923: inv_x_count_next = 16'b0000000001000111; // 1/923 = 0.0010834236
//      10'd924: inv_x_count_next = 16'b0000000001000111; // 1/924 = 0.0010822511
//      10'd925: inv_x_count_next = 16'b0000000001000111; // 1/925 = 0.0010810811
//      10'd926: inv_x_count_next = 16'b0000000001000111; // 1/926 = 0.0010799136
//      10'd927: inv_x_count_next = 16'b0000000001000111; // 1/927 = 0.0010787487
//      10'd928: inv_x_count_next = 16'b0000000001000111; // 1/928 = 0.0010775862
//      10'd929: inv_x_count_next = 16'b0000000001000111; // 1/929 = 0.0010764263
//      10'd930: inv_x_count_next = 16'b0000000001000110; // 1/930 = 0.0010752688
//      10'd931: inv_x_count_next = 16'b0000000001000110; // 1/931 = 0.0010741139
//      10'd932: inv_x_count_next = 16'b0000000001000110; // 1/932 = 0.0010729614
//      10'd933: inv_x_count_next = 16'b0000000001000110; // 1/933 = 0.0010718114
//      10'd934: inv_x_count_next = 16'b0000000001000110; // 1/934 = 0.0010706638
//      10'd935: inv_x_count_next = 16'b0000000001000110; // 1/935 = 0.0010695187
//      10'd936: inv_x_count_next = 16'b0000000001000110; // 1/936 = 0.0010683761
//      10'd937: inv_x_count_next = 16'b0000000001000110; // 1/937 = 0.0010672359
//      10'd938: inv_x_count_next = 16'b0000000001000110; // 1/938 = 0.0010660981
//      10'd939: inv_x_count_next = 16'b0000000001000110; // 1/939 = 0.0010649627
//      10'd940: inv_x_count_next = 16'b0000000001000110; // 1/940 = 0.0010638298
//      10'd941: inv_x_count_next = 16'b0000000001000110; // 1/941 = 0.0010626993
//      10'd942: inv_x_count_next = 16'b0000000001000110; // 1/942 = 0.0010615711
//      10'd943: inv_x_count_next = 16'b0000000001000101; // 1/943 = 0.0010604454
//      10'd944: inv_x_count_next = 16'b0000000001000101; // 1/944 = 0.0010593220
//      10'd945: inv_x_count_next = 16'b0000000001000101; // 1/945 = 0.0010582011
//      10'd946: inv_x_count_next = 16'b0000000001000101; // 1/946 = 0.0010570825
//      10'd947: inv_x_count_next = 16'b0000000001000101; // 1/947 = 0.0010559662
//      10'd948: inv_x_count_next = 16'b0000000001000101; // 1/948 = 0.0010548523
//      10'd949: inv_x_count_next = 16'b0000000001000101; // 1/949 = 0.0010537408
//      10'd950: inv_x_count_next = 16'b0000000001000101; // 1/950 = 0.0010526316
//      10'd951: inv_x_count_next = 16'b0000000001000101; // 1/951 = 0.0010515247
//      10'd952: inv_x_count_next = 16'b0000000001000101; // 1/952 = 0.0010504202
//      10'd953: inv_x_count_next = 16'b0000000001000101; // 1/953 = 0.0010493179
//      10'd954: inv_x_count_next = 16'b0000000001000101; // 1/954 = 0.0010482180
//      10'd955: inv_x_count_next = 16'b0000000001000101; // 1/955 = 0.0010471204
//      10'd956: inv_x_count_next = 16'b0000000001000101; // 1/956 = 0.0010460251
//      10'd957: inv_x_count_next = 16'b0000000001000100; // 1/957 = 0.0010449321
//      10'd958: inv_x_count_next = 16'b0000000001000100; // 1/958 = 0.0010438413
//      10'd959: inv_x_count_next = 16'b0000000001000100; // 1/959 = 0.0010427529
//      10'd960: inv_x_count_next = 16'b0000000001000100; // 1/960 = 0.0010416667
//      10'd961: inv_x_count_next = 16'b0000000001000100; // 1/961 = 0.0010405827
//      10'd962: inv_x_count_next = 16'b0000000001000100; // 1/962 = 0.0010395010
//      10'd963: inv_x_count_next = 16'b0000000001000100; // 1/963 = 0.0010384216
//      10'd964: inv_x_count_next = 16'b0000000001000100; // 1/964 = 0.0010373444
//      10'd965: inv_x_count_next = 16'b0000000001000100; // 1/965 = 0.0010362694
//      10'd966: inv_x_count_next = 16'b0000000001000100; // 1/966 = 0.0010351967
//      10'd967: inv_x_count_next = 16'b0000000001000100; // 1/967 = 0.0010341262
//      10'd968: inv_x_count_next = 16'b0000000001000100; // 1/968 = 0.0010330579
//      10'd969: inv_x_count_next = 16'b0000000001000100; // 1/969 = 0.0010319917
//      10'd970: inv_x_count_next = 16'b0000000001000100; // 1/970 = 0.0010309278
//      10'd971: inv_x_count_next = 16'b0000000001000011; // 1/971 = 0.0010298661
//      10'd972: inv_x_count_next = 16'b0000000001000011; // 1/972 = 0.0010288066
//      10'd973: inv_x_count_next = 16'b0000000001000011; // 1/973 = 0.0010277492
//      10'd974: inv_x_count_next = 16'b0000000001000011; // 1/974 = 0.0010266940
//      10'd975: inv_x_count_next = 16'b0000000001000011; // 1/975 = 0.0010256410
//      10'd976: inv_x_count_next = 16'b0000000001000011; // 1/976 = 0.0010245902
//      10'd977: inv_x_count_next = 16'b0000000001000011; // 1/977 = 0.0010235415
//      10'd978: inv_x_count_next = 16'b0000000001000011; // 1/978 = 0.0010224949
//      10'd979: inv_x_count_next = 16'b0000000001000011; // 1/979 = 0.0010214505
//      10'd980: inv_x_count_next = 16'b0000000001000011; // 1/980 = 0.0010204082
//      10'd981: inv_x_count_next = 16'b0000000001000011; // 1/981 = 0.0010193680
//      10'd982: inv_x_count_next = 16'b0000000001000011; // 1/982 = 0.0010183299
//      10'd983: inv_x_count_next = 16'b0000000001000011; // 1/983 = 0.0010172940
//      10'd984: inv_x_count_next = 16'b0000000001000011; // 1/984 = 0.0010162602
//      10'd985: inv_x_count_next = 16'b0000000001000011; // 1/985 = 0.0010152284
//      10'd986: inv_x_count_next = 16'b0000000001000010; // 1/986 = 0.0010141988
//      10'd987: inv_x_count_next = 16'b0000000001000010; // 1/987 = 0.0010131712
//      10'd988: inv_x_count_next = 16'b0000000001000010; // 1/988 = 0.0010121457
//      10'd989: inv_x_count_next = 16'b0000000001000010; // 1/989 = 0.0010111223
//      10'd990: inv_x_count_next = 16'b0000000001000010; // 1/990 = 0.0010101010
//      10'd991: inv_x_count_next = 16'b0000000001000010; // 1/991 = 0.0010090817
//      10'd992: inv_x_count_next = 16'b0000000001000010; // 1/992 = 0.0010080645
//      10'd993: inv_x_count_next = 16'b0000000001000010; // 1/993 = 0.0010070493
//      10'd994: inv_x_count_next = 16'b0000000001000010; // 1/994 = 0.0010060362
//      10'd995: inv_x_count_next = 16'b0000000001000010; // 1/995 = 0.0010050251
//      10'd996: inv_x_count_next = 16'b0000000001000010; // 1/996 = 0.0010040161
//      10'd997: inv_x_count_next = 16'b0000000001000010; // 1/997 = 0.0010030090
//      10'd998: inv_x_count_next = 16'b0000000001000010; // 1/998 = 0.0010020040
//      10'd999: inv_x_count_next = 16'b0000000001000010; // 1/999 = 0.0010010010
//      10'd1000: inv_x_count_next = 16'b0000000001000010; // 1/1000 = 0.0010000000
//      10'd1001: inv_x_count_next = 16'b0000000001000001; // 1/1001 = 0.0009990010
//      10'd1002: inv_x_count_next = 16'b0000000001000001; // 1/1002 = 0.0009980040
//      10'd1003: inv_x_count_next = 16'b0000000001000001; // 1/1003 = 0.0009970090
//      10'd1004: inv_x_count_next = 16'b0000000001000001; // 1/1004 = 0.0009960159
//      10'd1005: inv_x_count_next = 16'b0000000001000001; // 1/1005 = 0.0009950249
//      10'd1006: inv_x_count_next = 16'b0000000001000001; // 1/1006 = 0.0009940358
//      10'd1007: inv_x_count_next = 16'b0000000001000001; // 1/1007 = 0.0009930487
//      10'd1008: inv_x_count_next = 16'b0000000001000001; // 1/1008 = 0.0009920635
//      10'd1009: inv_x_count_next = 16'b0000000001000001; // 1/1009 = 0.0009910803
//      10'd1010: inv_x_count_next = 16'b0000000001000001; // 1/1010 = 0.0009900990
//      10'd1011: inv_x_count_next = 16'b0000000001000001; // 1/1011 = 0.0009891197
//      10'd1012: inv_x_count_next = 16'b0000000001000001; // 1/1012 = 0.0009881423
//      10'd1013: inv_x_count_next = 16'b0000000001000001; // 1/1013 = 0.0009871668
//      10'd1014: inv_x_count_next = 16'b0000000001000001; // 1/1014 = 0.0009861933
//      10'd1015: inv_x_count_next = 16'b0000000001000001; // 1/1015 = 0.0009852217
//      10'd1016: inv_x_count_next = 16'b0000000001000001; // 1/1016 = 0.0009842520
//      10'd1017: inv_x_count_next = 16'b0000000001000000; // 1/1017 = 0.0009832842
//      10'd1018: inv_x_count_next = 16'b0000000001000000; // 1/1018 = 0.0009823183
//      10'd1019: inv_x_count_next = 16'b0000000001000000; // 1/1019 = 0.0009813543
//      10'd1020: inv_x_count_next = 16'b0000000001000000; // 1/1020 = 0.0009803922
//      10'd1021: inv_x_count_next = 16'b0000000001000000; // 1/1021 = 0.0009794319
//      10'd1022: inv_x_count_next = 16'b0000000001000000; // 1/1022 = 0.0009784736
//      10'd1023: inv_x_count_next = 16'b0000000001000000; // 1/1023 = 0.0009775171
//      10'd1024: inv_x_count_next = 16'b0000000001000000; // 1/1024 = 0.0009765625
//      default: inv_x_count_next = '0; // Default case
//    endcase
//  end
endmodule
